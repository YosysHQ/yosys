// Created by cells_xtra.py from Xilinx models

module CMAC (...);
    parameter CTL_PTP_TRANSPCLK_MODE = "FALSE";
    parameter CTL_RX_CHECK_ACK = "TRUE";
    parameter CTL_RX_CHECK_PREAMBLE = "FALSE";
    parameter CTL_RX_CHECK_SFD = "FALSE";
    parameter CTL_RX_DELETE_FCS = "TRUE";
    parameter [15:0] CTL_RX_ETYPE_GCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_GPP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PPP = 16'h8808;
    parameter CTL_RX_FORWARD_CONTROL = "FALSE";
    parameter CTL_RX_IGNORE_FCS = "FALSE";
    parameter [14:0] CTL_RX_MAX_PACKET_LEN = 15'h2580;
    parameter [7:0] CTL_RX_MIN_PACKET_LEN = 8'h40;
    parameter [15:0] CTL_RX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_RX_OPCODE_MAX_GCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MAX_PCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MIN_GCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_MIN_PCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_PPP = 16'h0001;
    parameter [47:0] CTL_RX_PAUSE_DA_MCAST = 48'h0180C2000001;
    parameter [47:0] CTL_RX_PAUSE_DA_UCAST = 48'h000000000000;
    parameter [47:0] CTL_RX_PAUSE_SA = 48'h000000000000;
    parameter CTL_RX_PROCESS_LFI = "FALSE";
    parameter [15:0] CTL_RX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_RX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_RX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_RX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_RX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_RX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_RX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_RX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_RX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_RX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_RX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_RX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_RX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_RX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_RX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_RX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_RX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_RX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_RX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [47:0] CTL_TX_DA_GPP = 48'h0180C2000001;
    parameter [47:0] CTL_TX_DA_PPP = 48'h0180C2000001;
    parameter [15:0] CTL_TX_ETHERTYPE_GPP = 16'h8808;
    parameter [15:0] CTL_TX_ETHERTYPE_PPP = 16'h8808;
    parameter CTL_TX_FCS_INS_ENABLE = "TRUE";
    parameter CTL_TX_IGNORE_FCS = "FALSE";
    parameter [15:0] CTL_TX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_TX_OPCODE_PPP = 16'h0001;
    parameter CTL_TX_PTP_1STEP_ENABLE = "FALSE";
    parameter [10:0] CTL_TX_PTP_LATENCY_ADJUST = 11'h2C1;
    parameter [47:0] CTL_TX_SA_GPP = 48'h000000000000;
    parameter [47:0] CTL_TX_SA_PPP = 48'h000000000000;
    parameter [15:0] CTL_TX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_TX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_TX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_TX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_TX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_TX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_TX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_TX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_TX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_TX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_TX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_TX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_TX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_TX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_TX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_TX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_TX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_TX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_TX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter SIM_VERSION = "2.0";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [6:0] RX_LANE_ALIGNER_FILL_0;
    output [6:0] RX_LANE_ALIGNER_FILL_1;
    output [6:0] RX_LANE_ALIGNER_FILL_10;
    output [6:0] RX_LANE_ALIGNER_FILL_11;
    output [6:0] RX_LANE_ALIGNER_FILL_12;
    output [6:0] RX_LANE_ALIGNER_FILL_13;
    output [6:0] RX_LANE_ALIGNER_FILL_14;
    output [6:0] RX_LANE_ALIGNER_FILL_15;
    output [6:0] RX_LANE_ALIGNER_FILL_16;
    output [6:0] RX_LANE_ALIGNER_FILL_17;
    output [6:0] RX_LANE_ALIGNER_FILL_18;
    output [6:0] RX_LANE_ALIGNER_FILL_19;
    output [6:0] RX_LANE_ALIGNER_FILL_2;
    output [6:0] RX_LANE_ALIGNER_FILL_3;
    output [6:0] RX_LANE_ALIGNER_FILL_4;
    output [6:0] RX_LANE_ALIGNER_FILL_5;
    output [6:0] RX_LANE_ALIGNER_FILL_6;
    output [6:0] RX_LANE_ALIGNER_FILL_7;
    output [6:0] RX_LANE_ALIGNER_FILL_8;
    output [6:0] RX_LANE_ALIGNER_FILL_9;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output [4:0] RX_PTP_PCSLANE_OUT;
    output [79:0] RX_PTP_TSTAMP_OUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [6:0] STAT_RX_BAD_CODE;
    output [3:0] STAT_RX_BAD_FCS;
    output STAT_RX_BAD_PREAMBLE;
    output STAT_RX_BAD_SFD;
    output STAT_RX_BIP_ERR_0;
    output STAT_RX_BIP_ERR_1;
    output STAT_RX_BIP_ERR_10;
    output STAT_RX_BIP_ERR_11;
    output STAT_RX_BIP_ERR_12;
    output STAT_RX_BIP_ERR_13;
    output STAT_RX_BIP_ERR_14;
    output STAT_RX_BIP_ERR_15;
    output STAT_RX_BIP_ERR_16;
    output STAT_RX_BIP_ERR_17;
    output STAT_RX_BIP_ERR_18;
    output STAT_RX_BIP_ERR_19;
    output STAT_RX_BIP_ERR_2;
    output STAT_RX_BIP_ERR_3;
    output STAT_RX_BIP_ERR_4;
    output STAT_RX_BIP_ERR_5;
    output STAT_RX_BIP_ERR_6;
    output STAT_RX_BIP_ERR_7;
    output STAT_RX_BIP_ERR_8;
    output STAT_RX_BIP_ERR_9;
    output [19:0] STAT_RX_BLOCK_LOCK;
    output STAT_RX_BROADCAST;
    output [3:0] STAT_RX_FRAGMENT;
    output [3:0] STAT_RX_FRAMING_ERR_0;
    output [3:0] STAT_RX_FRAMING_ERR_1;
    output [3:0] STAT_RX_FRAMING_ERR_10;
    output [3:0] STAT_RX_FRAMING_ERR_11;
    output [3:0] STAT_RX_FRAMING_ERR_12;
    output [3:0] STAT_RX_FRAMING_ERR_13;
    output [3:0] STAT_RX_FRAMING_ERR_14;
    output [3:0] STAT_RX_FRAMING_ERR_15;
    output [3:0] STAT_RX_FRAMING_ERR_16;
    output [3:0] STAT_RX_FRAMING_ERR_17;
    output [3:0] STAT_RX_FRAMING_ERR_18;
    output [3:0] STAT_RX_FRAMING_ERR_19;
    output [3:0] STAT_RX_FRAMING_ERR_2;
    output [3:0] STAT_RX_FRAMING_ERR_3;
    output [3:0] STAT_RX_FRAMING_ERR_4;
    output [3:0] STAT_RX_FRAMING_ERR_5;
    output [3:0] STAT_RX_FRAMING_ERR_6;
    output [3:0] STAT_RX_FRAMING_ERR_7;
    output [3:0] STAT_RX_FRAMING_ERR_8;
    output [3:0] STAT_RX_FRAMING_ERR_9;
    output STAT_RX_FRAMING_ERR_VALID_0;
    output STAT_RX_FRAMING_ERR_VALID_1;
    output STAT_RX_FRAMING_ERR_VALID_10;
    output STAT_RX_FRAMING_ERR_VALID_11;
    output STAT_RX_FRAMING_ERR_VALID_12;
    output STAT_RX_FRAMING_ERR_VALID_13;
    output STAT_RX_FRAMING_ERR_VALID_14;
    output STAT_RX_FRAMING_ERR_VALID_15;
    output STAT_RX_FRAMING_ERR_VALID_16;
    output STAT_RX_FRAMING_ERR_VALID_17;
    output STAT_RX_FRAMING_ERR_VALID_18;
    output STAT_RX_FRAMING_ERR_VALID_19;
    output STAT_RX_FRAMING_ERR_VALID_2;
    output STAT_RX_FRAMING_ERR_VALID_3;
    output STAT_RX_FRAMING_ERR_VALID_4;
    output STAT_RX_FRAMING_ERR_VALID_5;
    output STAT_RX_FRAMING_ERR_VALID_6;
    output STAT_RX_FRAMING_ERR_VALID_7;
    output STAT_RX_FRAMING_ERR_VALID_8;
    output STAT_RX_FRAMING_ERR_VALID_9;
    output STAT_RX_GOT_SIGNAL_OS;
    output STAT_RX_HI_BER;
    output STAT_RX_INRANGEERR;
    output STAT_RX_INTERNAL_LOCAL_FAULT;
    output STAT_RX_JABBER;
    output [7:0] STAT_RX_LANE0_VLM_BIP7;
    output STAT_RX_LANE0_VLM_BIP7_VALID;
    output STAT_RX_LOCAL_FAULT;
    output [19:0] STAT_RX_MF_ERR;
    output [19:0] STAT_RX_MF_LEN_ERR;
    output [19:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MULTICAST;
    output STAT_RX_OVERSIZE;
    output STAT_RX_PACKET_1024_1518_BYTES;
    output STAT_RX_PACKET_128_255_BYTES;
    output STAT_RX_PACKET_1519_1522_BYTES;
    output STAT_RX_PACKET_1523_1548_BYTES;
    output STAT_RX_PACKET_1549_2047_BYTES;
    output STAT_RX_PACKET_2048_4095_BYTES;
    output STAT_RX_PACKET_256_511_BYTES;
    output STAT_RX_PACKET_4096_8191_BYTES;
    output STAT_RX_PACKET_512_1023_BYTES;
    output STAT_RX_PACKET_64_BYTES;
    output STAT_RX_PACKET_65_127_BYTES;
    output STAT_RX_PACKET_8192_9215_BYTES;
    output STAT_RX_PACKET_BAD_FCS;
    output STAT_RX_PACKET_LARGE;
    output [3:0] STAT_RX_PACKET_SMALL;
    output STAT_RX_PAUSE;
    output [15:0] STAT_RX_PAUSE_QUANTA0;
    output [15:0] STAT_RX_PAUSE_QUANTA1;
    output [15:0] STAT_RX_PAUSE_QUANTA2;
    output [15:0] STAT_RX_PAUSE_QUANTA3;
    output [15:0] STAT_RX_PAUSE_QUANTA4;
    output [15:0] STAT_RX_PAUSE_QUANTA5;
    output [15:0] STAT_RX_PAUSE_QUANTA6;
    output [15:0] STAT_RX_PAUSE_QUANTA7;
    output [15:0] STAT_RX_PAUSE_QUANTA8;
    output [8:0] STAT_RX_PAUSE_REQ;
    output [8:0] STAT_RX_PAUSE_VALID;
    output STAT_RX_RECEIVED_LOCAL_FAULT;
    output STAT_RX_REMOTE_FAULT;
    output STAT_RX_STATUS;
    output [3:0] STAT_RX_STOMPED_FCS;
    output [19:0] STAT_RX_SYNCED;
    output [19:0] STAT_RX_SYNCED_ERR;
    output [2:0] STAT_RX_TEST_PATTERN_MISMATCH;
    output STAT_RX_TOOLONG;
    output [7:0] STAT_RX_TOTAL_BYTES;
    output [13:0] STAT_RX_TOTAL_GOOD_BYTES;
    output STAT_RX_TOTAL_GOOD_PACKETS;
    output [3:0] STAT_RX_TOTAL_PACKETS;
    output STAT_RX_TRUNCATED;
    output [3:0] STAT_RX_UNDERSIZE;
    output STAT_RX_UNICAST;
    output STAT_RX_USER_PAUSE;
    output STAT_RX_VLAN;
    output [19:0] STAT_RX_VL_DEMUXED;
    output [4:0] STAT_RX_VL_NUMBER_0;
    output [4:0] STAT_RX_VL_NUMBER_1;
    output [4:0] STAT_RX_VL_NUMBER_10;
    output [4:0] STAT_RX_VL_NUMBER_11;
    output [4:0] STAT_RX_VL_NUMBER_12;
    output [4:0] STAT_RX_VL_NUMBER_13;
    output [4:0] STAT_RX_VL_NUMBER_14;
    output [4:0] STAT_RX_VL_NUMBER_15;
    output [4:0] STAT_RX_VL_NUMBER_16;
    output [4:0] STAT_RX_VL_NUMBER_17;
    output [4:0] STAT_RX_VL_NUMBER_18;
    output [4:0] STAT_RX_VL_NUMBER_19;
    output [4:0] STAT_RX_VL_NUMBER_2;
    output [4:0] STAT_RX_VL_NUMBER_3;
    output [4:0] STAT_RX_VL_NUMBER_4;
    output [4:0] STAT_RX_VL_NUMBER_5;
    output [4:0] STAT_RX_VL_NUMBER_6;
    output [4:0] STAT_RX_VL_NUMBER_7;
    output [4:0] STAT_RX_VL_NUMBER_8;
    output [4:0] STAT_RX_VL_NUMBER_9;
    output STAT_TX_BAD_FCS;
    output STAT_TX_BROADCAST;
    output STAT_TX_FRAME_ERROR;
    output STAT_TX_LOCAL_FAULT;
    output STAT_TX_MULTICAST;
    output STAT_TX_PACKET_1024_1518_BYTES;
    output STAT_TX_PACKET_128_255_BYTES;
    output STAT_TX_PACKET_1519_1522_BYTES;
    output STAT_TX_PACKET_1523_1548_BYTES;
    output STAT_TX_PACKET_1549_2047_BYTES;
    output STAT_TX_PACKET_2048_4095_BYTES;
    output STAT_TX_PACKET_256_511_BYTES;
    output STAT_TX_PACKET_4096_8191_BYTES;
    output STAT_TX_PACKET_512_1023_BYTES;
    output STAT_TX_PACKET_64_BYTES;
    output STAT_TX_PACKET_65_127_BYTES;
    output STAT_TX_PACKET_8192_9215_BYTES;
    output STAT_TX_PACKET_LARGE;
    output STAT_TX_PACKET_SMALL;
    output STAT_TX_PAUSE;
    output [8:0] STAT_TX_PAUSE_VALID;
    output STAT_TX_PTP_FIFO_READ_ERROR;
    output STAT_TX_PTP_FIFO_WRITE_ERROR;
    output [6:0] STAT_TX_TOTAL_BYTES;
    output [13:0] STAT_TX_TOTAL_GOOD_BYTES;
    output STAT_TX_TOTAL_GOOD_PACKETS;
    output STAT_TX_TOTAL_PACKETS;
    output STAT_TX_UNICAST;
    output STAT_TX_USER_PAUSE;
    output STAT_TX_VLAN;
    output TX_OVFOUT;
    output [4:0] TX_PTP_PCSLANE_OUT;
    output [79:0] TX_PTP_TSTAMP_OUT;
    output [15:0] TX_PTP_TSTAMP_TAG_OUT;
    output TX_PTP_TSTAMP_VALID_OUT;
    output TX_RDYOUT;
    output [15:0] TX_SERDES_ALT_DATA0;
    output [15:0] TX_SERDES_ALT_DATA1;
    output [15:0] TX_SERDES_ALT_DATA2;
    output [15:0] TX_SERDES_ALT_DATA3;
    output [63:0] TX_SERDES_DATA0;
    output [63:0] TX_SERDES_DATA1;
    output [63:0] TX_SERDES_DATA2;
    output [63:0] TX_SERDES_DATA3;
    output [31:0] TX_SERDES_DATA4;
    output [31:0] TX_SERDES_DATA5;
    output [31:0] TX_SERDES_DATA6;
    output [31:0] TX_SERDES_DATA7;
    output [31:0] TX_SERDES_DATA8;
    output [31:0] TX_SERDES_DATA9;
    output TX_UNFOUT;
    input CTL_CAUI4_MODE;
    input CTL_RX_CHECK_ETYPE_GCP;
    input CTL_RX_CHECK_ETYPE_GPP;
    input CTL_RX_CHECK_ETYPE_PCP;
    input CTL_RX_CHECK_ETYPE_PPP;
    input CTL_RX_CHECK_MCAST_GCP;
    input CTL_RX_CHECK_MCAST_GPP;
    input CTL_RX_CHECK_MCAST_PCP;
    input CTL_RX_CHECK_MCAST_PPP;
    input CTL_RX_CHECK_OPCODE_GCP;
    input CTL_RX_CHECK_OPCODE_GPP;
    input CTL_RX_CHECK_OPCODE_PCP;
    input CTL_RX_CHECK_OPCODE_PPP;
    input CTL_RX_CHECK_SA_GCP;
    input CTL_RX_CHECK_SA_GPP;
    input CTL_RX_CHECK_SA_PCP;
    input CTL_RX_CHECK_SA_PPP;
    input CTL_RX_CHECK_UCAST_GCP;
    input CTL_RX_CHECK_UCAST_GPP;
    input CTL_RX_CHECK_UCAST_PCP;
    input CTL_RX_CHECK_UCAST_PPP;
    input CTL_RX_ENABLE;
    input CTL_RX_ENABLE_GCP;
    input CTL_RX_ENABLE_GPP;
    input CTL_RX_ENABLE_PCP;
    input CTL_RX_ENABLE_PPP;
    input CTL_RX_FORCE_RESYNC;
    input [8:0] CTL_RX_PAUSE_ACK;
    input [8:0] CTL_RX_PAUSE_ENABLE;
    input [79:0] CTL_RX_SYSTEMTIMERIN;
    input CTL_RX_TEST_PATTERN;
    input CTL_TX_ENABLE;
    input CTL_TX_LANE0_VLM_BIP7_OVERRIDE;
    input [7:0] CTL_TX_LANE0_VLM_BIP7_OVERRIDE_VALUE;
    input [8:0] CTL_TX_PAUSE_ENABLE;
    input [15:0] CTL_TX_PAUSE_QUANTA0;
    input [15:0] CTL_TX_PAUSE_QUANTA1;
    input [15:0] CTL_TX_PAUSE_QUANTA2;
    input [15:0] CTL_TX_PAUSE_QUANTA3;
    input [15:0] CTL_TX_PAUSE_QUANTA4;
    input [15:0] CTL_TX_PAUSE_QUANTA5;
    input [15:0] CTL_TX_PAUSE_QUANTA6;
    input [15:0] CTL_TX_PAUSE_QUANTA7;
    input [15:0] CTL_TX_PAUSE_QUANTA8;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER0;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER1;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER2;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER3;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER4;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER5;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER6;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER7;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER8;
    input [8:0] CTL_TX_PAUSE_REQ;
    input CTL_TX_PTP_VLANE_ADJUST_MODE;
    input CTL_TX_RESEND_PAUSE;
    input CTL_TX_SEND_IDLE;
    input CTL_TX_SEND_RFI;
    input [79:0] CTL_TX_SYSTEMTIMERIN;
    input CTL_TX_TEST_PATTERN;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input RX_CLK;
    input RX_RESET;
    input [15:0] RX_SERDES_ALT_DATA0;
    input [15:0] RX_SERDES_ALT_DATA1;
    input [15:0] RX_SERDES_ALT_DATA2;
    input [15:0] RX_SERDES_ALT_DATA3;
    input [9:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA0;
    input [63:0] RX_SERDES_DATA1;
    input [63:0] RX_SERDES_DATA2;
    input [63:0] RX_SERDES_DATA3;
    input [31:0] RX_SERDES_DATA4;
    input [31:0] RX_SERDES_DATA5;
    input [31:0] RX_SERDES_DATA6;
    input [31:0] RX_SERDES_DATA7;
    input [31:0] RX_SERDES_DATA8;
    input [31:0] RX_SERDES_DATA9;
    input [9:0] RX_SERDES_RESET;
    input TX_CLK;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input [1:0] TX_PTP_1588OP_IN;
    input [15:0] TX_PTP_CHKSUM_OFFSET_IN;
    input [63:0] TX_PTP_RXTSTAMP_IN;
    input [15:0] TX_PTP_TAG_FIELD_IN;
    input [15:0] TX_PTP_TSTAMP_OFFSET_IN;
    input TX_PTP_UPD_CHKSUM_IN;
    input TX_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module CMACE4 (...);
    parameter CTL_PTP_TRANSPCLK_MODE = "FALSE";
    parameter CTL_RX_CHECK_ACK = "TRUE";
    parameter CTL_RX_CHECK_PREAMBLE = "FALSE";
    parameter CTL_RX_CHECK_SFD = "FALSE";
    parameter CTL_RX_DELETE_FCS = "TRUE";
    parameter [15:0] CTL_RX_ETYPE_GCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_GPP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PPP = 16'h8808;
    parameter CTL_RX_FORWARD_CONTROL = "FALSE";
    parameter CTL_RX_IGNORE_FCS = "FALSE";
    parameter [14:0] CTL_RX_MAX_PACKET_LEN = 15'h2580;
    parameter [7:0] CTL_RX_MIN_PACKET_LEN = 8'h40;
    parameter [15:0] CTL_RX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_RX_OPCODE_MAX_GCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MAX_PCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MIN_GCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_MIN_PCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_PPP = 16'h0001;
    parameter [47:0] CTL_RX_PAUSE_DA_MCAST = 48'h0180C2000001;
    parameter [47:0] CTL_RX_PAUSE_DA_UCAST = 48'h000000000000;
    parameter [47:0] CTL_RX_PAUSE_SA = 48'h000000000000;
    parameter CTL_RX_PROCESS_LFI = "FALSE";
    parameter [8:0] CTL_RX_RSFEC_AM_THRESHOLD = 9'h046;
    parameter [1:0] CTL_RX_RSFEC_FILL_ADJUST = 2'h0;
    parameter [15:0] CTL_RX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_RX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_RX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_RX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_RX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_RX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_RX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_RX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_RX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_RX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_RX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_RX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_RX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_RX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_RX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_RX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_RX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_RX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_RX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter CTL_TX_CUSTOM_PREAMBLE_ENABLE = "FALSE";
    parameter [47:0] CTL_TX_DA_GPP = 48'h0180C2000001;
    parameter [47:0] CTL_TX_DA_PPP = 48'h0180C2000001;
    parameter [15:0] CTL_TX_ETHERTYPE_GPP = 16'h8808;
    parameter [15:0] CTL_TX_ETHERTYPE_PPP = 16'h8808;
    parameter CTL_TX_FCS_INS_ENABLE = "TRUE";
    parameter CTL_TX_IGNORE_FCS = "FALSE";
    parameter [3:0] CTL_TX_IPG_VALUE = 4'hC;
    parameter [15:0] CTL_TX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_TX_OPCODE_PPP = 16'h0001;
    parameter CTL_TX_PTP_1STEP_ENABLE = "FALSE";
    parameter [10:0] CTL_TX_PTP_LATENCY_ADJUST = 11'h2C1;
    parameter [47:0] CTL_TX_SA_GPP = 48'h000000000000;
    parameter [47:0] CTL_TX_SA_PPP = 48'h000000000000;
    parameter [15:0] CTL_TX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_TX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_TX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_TX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_TX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_TX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_TX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_TX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_TX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_TX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_TX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_TX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_TX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_TX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_TX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_TX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_TX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_TX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_TX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [329:0] RSFEC_BYPASS_RX_DOUT;
    output RSFEC_BYPASS_RX_DOUT_CW_START;
    output RSFEC_BYPASS_RX_DOUT_VALID;
    output [329:0] RSFEC_BYPASS_TX_DOUT;
    output RSFEC_BYPASS_TX_DOUT_CW_START;
    output RSFEC_BYPASS_TX_DOUT_VALID;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [6:0] RX_LANE_ALIGNER_FILL_0;
    output [6:0] RX_LANE_ALIGNER_FILL_1;
    output [6:0] RX_LANE_ALIGNER_FILL_10;
    output [6:0] RX_LANE_ALIGNER_FILL_11;
    output [6:0] RX_LANE_ALIGNER_FILL_12;
    output [6:0] RX_LANE_ALIGNER_FILL_13;
    output [6:0] RX_LANE_ALIGNER_FILL_14;
    output [6:0] RX_LANE_ALIGNER_FILL_15;
    output [6:0] RX_LANE_ALIGNER_FILL_16;
    output [6:0] RX_LANE_ALIGNER_FILL_17;
    output [6:0] RX_LANE_ALIGNER_FILL_18;
    output [6:0] RX_LANE_ALIGNER_FILL_19;
    output [6:0] RX_LANE_ALIGNER_FILL_2;
    output [6:0] RX_LANE_ALIGNER_FILL_3;
    output [6:0] RX_LANE_ALIGNER_FILL_4;
    output [6:0] RX_LANE_ALIGNER_FILL_5;
    output [6:0] RX_LANE_ALIGNER_FILL_6;
    output [6:0] RX_LANE_ALIGNER_FILL_7;
    output [6:0] RX_LANE_ALIGNER_FILL_8;
    output [6:0] RX_LANE_ALIGNER_FILL_9;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output [7:0] RX_OTN_BIP8_0;
    output [7:0] RX_OTN_BIP8_1;
    output [7:0] RX_OTN_BIP8_2;
    output [7:0] RX_OTN_BIP8_3;
    output [7:0] RX_OTN_BIP8_4;
    output [65:0] RX_OTN_DATA_0;
    output [65:0] RX_OTN_DATA_1;
    output [65:0] RX_OTN_DATA_2;
    output [65:0] RX_OTN_DATA_3;
    output [65:0] RX_OTN_DATA_4;
    output RX_OTN_ENA;
    output RX_OTN_LANE0;
    output RX_OTN_VLMARKER;
    output [55:0] RX_PREOUT;
    output [4:0] RX_PTP_PCSLANE_OUT;
    output [79:0] RX_PTP_TSTAMP_OUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [2:0] STAT_RX_BAD_CODE;
    output [2:0] STAT_RX_BAD_FCS;
    output STAT_RX_BAD_PREAMBLE;
    output STAT_RX_BAD_SFD;
    output STAT_RX_BIP_ERR_0;
    output STAT_RX_BIP_ERR_1;
    output STAT_RX_BIP_ERR_10;
    output STAT_RX_BIP_ERR_11;
    output STAT_RX_BIP_ERR_12;
    output STAT_RX_BIP_ERR_13;
    output STAT_RX_BIP_ERR_14;
    output STAT_RX_BIP_ERR_15;
    output STAT_RX_BIP_ERR_16;
    output STAT_RX_BIP_ERR_17;
    output STAT_RX_BIP_ERR_18;
    output STAT_RX_BIP_ERR_19;
    output STAT_RX_BIP_ERR_2;
    output STAT_RX_BIP_ERR_3;
    output STAT_RX_BIP_ERR_4;
    output STAT_RX_BIP_ERR_5;
    output STAT_RX_BIP_ERR_6;
    output STAT_RX_BIP_ERR_7;
    output STAT_RX_BIP_ERR_8;
    output STAT_RX_BIP_ERR_9;
    output [19:0] STAT_RX_BLOCK_LOCK;
    output STAT_RX_BROADCAST;
    output [2:0] STAT_RX_FRAGMENT;
    output [1:0] STAT_RX_FRAMING_ERR_0;
    output [1:0] STAT_RX_FRAMING_ERR_1;
    output [1:0] STAT_RX_FRAMING_ERR_10;
    output [1:0] STAT_RX_FRAMING_ERR_11;
    output [1:0] STAT_RX_FRAMING_ERR_12;
    output [1:0] STAT_RX_FRAMING_ERR_13;
    output [1:0] STAT_RX_FRAMING_ERR_14;
    output [1:0] STAT_RX_FRAMING_ERR_15;
    output [1:0] STAT_RX_FRAMING_ERR_16;
    output [1:0] STAT_RX_FRAMING_ERR_17;
    output [1:0] STAT_RX_FRAMING_ERR_18;
    output [1:0] STAT_RX_FRAMING_ERR_19;
    output [1:0] STAT_RX_FRAMING_ERR_2;
    output [1:0] STAT_RX_FRAMING_ERR_3;
    output [1:0] STAT_RX_FRAMING_ERR_4;
    output [1:0] STAT_RX_FRAMING_ERR_5;
    output [1:0] STAT_RX_FRAMING_ERR_6;
    output [1:0] STAT_RX_FRAMING_ERR_7;
    output [1:0] STAT_RX_FRAMING_ERR_8;
    output [1:0] STAT_RX_FRAMING_ERR_9;
    output STAT_RX_FRAMING_ERR_VALID_0;
    output STAT_RX_FRAMING_ERR_VALID_1;
    output STAT_RX_FRAMING_ERR_VALID_10;
    output STAT_RX_FRAMING_ERR_VALID_11;
    output STAT_RX_FRAMING_ERR_VALID_12;
    output STAT_RX_FRAMING_ERR_VALID_13;
    output STAT_RX_FRAMING_ERR_VALID_14;
    output STAT_RX_FRAMING_ERR_VALID_15;
    output STAT_RX_FRAMING_ERR_VALID_16;
    output STAT_RX_FRAMING_ERR_VALID_17;
    output STAT_RX_FRAMING_ERR_VALID_18;
    output STAT_RX_FRAMING_ERR_VALID_19;
    output STAT_RX_FRAMING_ERR_VALID_2;
    output STAT_RX_FRAMING_ERR_VALID_3;
    output STAT_RX_FRAMING_ERR_VALID_4;
    output STAT_RX_FRAMING_ERR_VALID_5;
    output STAT_RX_FRAMING_ERR_VALID_6;
    output STAT_RX_FRAMING_ERR_VALID_7;
    output STAT_RX_FRAMING_ERR_VALID_8;
    output STAT_RX_FRAMING_ERR_VALID_9;
    output STAT_RX_GOT_SIGNAL_OS;
    output STAT_RX_HI_BER;
    output STAT_RX_INRANGEERR;
    output STAT_RX_INTERNAL_LOCAL_FAULT;
    output STAT_RX_JABBER;
    output [7:0] STAT_RX_LANE0_VLM_BIP7;
    output STAT_RX_LANE0_VLM_BIP7_VALID;
    output STAT_RX_LOCAL_FAULT;
    output [19:0] STAT_RX_MF_ERR;
    output [19:0] STAT_RX_MF_LEN_ERR;
    output [19:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MULTICAST;
    output STAT_RX_OVERSIZE;
    output STAT_RX_PACKET_1024_1518_BYTES;
    output STAT_RX_PACKET_128_255_BYTES;
    output STAT_RX_PACKET_1519_1522_BYTES;
    output STAT_RX_PACKET_1523_1548_BYTES;
    output STAT_RX_PACKET_1549_2047_BYTES;
    output STAT_RX_PACKET_2048_4095_BYTES;
    output STAT_RX_PACKET_256_511_BYTES;
    output STAT_RX_PACKET_4096_8191_BYTES;
    output STAT_RX_PACKET_512_1023_BYTES;
    output STAT_RX_PACKET_64_BYTES;
    output STAT_RX_PACKET_65_127_BYTES;
    output STAT_RX_PACKET_8192_9215_BYTES;
    output STAT_RX_PACKET_BAD_FCS;
    output STAT_RX_PACKET_LARGE;
    output [2:0] STAT_RX_PACKET_SMALL;
    output STAT_RX_PAUSE;
    output [15:0] STAT_RX_PAUSE_QUANTA0;
    output [15:0] STAT_RX_PAUSE_QUANTA1;
    output [15:0] STAT_RX_PAUSE_QUANTA2;
    output [15:0] STAT_RX_PAUSE_QUANTA3;
    output [15:0] STAT_RX_PAUSE_QUANTA4;
    output [15:0] STAT_RX_PAUSE_QUANTA5;
    output [15:0] STAT_RX_PAUSE_QUANTA6;
    output [15:0] STAT_RX_PAUSE_QUANTA7;
    output [15:0] STAT_RX_PAUSE_QUANTA8;
    output [8:0] STAT_RX_PAUSE_REQ;
    output [8:0] STAT_RX_PAUSE_VALID;
    output STAT_RX_RECEIVED_LOCAL_FAULT;
    output STAT_RX_REMOTE_FAULT;
    output STAT_RX_RSFEC_AM_LOCK0;
    output STAT_RX_RSFEC_AM_LOCK1;
    output STAT_RX_RSFEC_AM_LOCK2;
    output STAT_RX_RSFEC_AM_LOCK3;
    output STAT_RX_RSFEC_CORRECTED_CW_INC;
    output STAT_RX_RSFEC_CW_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT0_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT1_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT2_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT3_INC;
    output STAT_RX_RSFEC_HI_SER;
    output STAT_RX_RSFEC_LANE_ALIGNMENT_STATUS;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_0;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_1;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_2;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_3;
    output [7:0] STAT_RX_RSFEC_LANE_MAPPING;
    output [31:0] STAT_RX_RSFEC_RSVD;
    output STAT_RX_RSFEC_UNCORRECTED_CW_INC;
    output STAT_RX_STATUS;
    output [2:0] STAT_RX_STOMPED_FCS;
    output [19:0] STAT_RX_SYNCED;
    output [19:0] STAT_RX_SYNCED_ERR;
    output [2:0] STAT_RX_TEST_PATTERN_MISMATCH;
    output STAT_RX_TOOLONG;
    output [6:0] STAT_RX_TOTAL_BYTES;
    output [13:0] STAT_RX_TOTAL_GOOD_BYTES;
    output STAT_RX_TOTAL_GOOD_PACKETS;
    output [2:0] STAT_RX_TOTAL_PACKETS;
    output STAT_RX_TRUNCATED;
    output [2:0] STAT_RX_UNDERSIZE;
    output STAT_RX_UNICAST;
    output STAT_RX_USER_PAUSE;
    output STAT_RX_VLAN;
    output [19:0] STAT_RX_VL_DEMUXED;
    output [4:0] STAT_RX_VL_NUMBER_0;
    output [4:0] STAT_RX_VL_NUMBER_1;
    output [4:0] STAT_RX_VL_NUMBER_10;
    output [4:0] STAT_RX_VL_NUMBER_11;
    output [4:0] STAT_RX_VL_NUMBER_12;
    output [4:0] STAT_RX_VL_NUMBER_13;
    output [4:0] STAT_RX_VL_NUMBER_14;
    output [4:0] STAT_RX_VL_NUMBER_15;
    output [4:0] STAT_RX_VL_NUMBER_16;
    output [4:0] STAT_RX_VL_NUMBER_17;
    output [4:0] STAT_RX_VL_NUMBER_18;
    output [4:0] STAT_RX_VL_NUMBER_19;
    output [4:0] STAT_RX_VL_NUMBER_2;
    output [4:0] STAT_RX_VL_NUMBER_3;
    output [4:0] STAT_RX_VL_NUMBER_4;
    output [4:0] STAT_RX_VL_NUMBER_5;
    output [4:0] STAT_RX_VL_NUMBER_6;
    output [4:0] STAT_RX_VL_NUMBER_7;
    output [4:0] STAT_RX_VL_NUMBER_8;
    output [4:0] STAT_RX_VL_NUMBER_9;
    output STAT_TX_BAD_FCS;
    output STAT_TX_BROADCAST;
    output STAT_TX_FRAME_ERROR;
    output STAT_TX_LOCAL_FAULT;
    output STAT_TX_MULTICAST;
    output STAT_TX_PACKET_1024_1518_BYTES;
    output STAT_TX_PACKET_128_255_BYTES;
    output STAT_TX_PACKET_1519_1522_BYTES;
    output STAT_TX_PACKET_1523_1548_BYTES;
    output STAT_TX_PACKET_1549_2047_BYTES;
    output STAT_TX_PACKET_2048_4095_BYTES;
    output STAT_TX_PACKET_256_511_BYTES;
    output STAT_TX_PACKET_4096_8191_BYTES;
    output STAT_TX_PACKET_512_1023_BYTES;
    output STAT_TX_PACKET_64_BYTES;
    output STAT_TX_PACKET_65_127_BYTES;
    output STAT_TX_PACKET_8192_9215_BYTES;
    output STAT_TX_PACKET_LARGE;
    output STAT_TX_PACKET_SMALL;
    output STAT_TX_PAUSE;
    output [8:0] STAT_TX_PAUSE_VALID;
    output STAT_TX_PTP_FIFO_READ_ERROR;
    output STAT_TX_PTP_FIFO_WRITE_ERROR;
    output [5:0] STAT_TX_TOTAL_BYTES;
    output [13:0] STAT_TX_TOTAL_GOOD_BYTES;
    output STAT_TX_TOTAL_GOOD_PACKETS;
    output STAT_TX_TOTAL_PACKETS;
    output STAT_TX_UNICAST;
    output STAT_TX_USER_PAUSE;
    output STAT_TX_VLAN;
    output TX_OVFOUT;
    output [4:0] TX_PTP_PCSLANE_OUT;
    output [79:0] TX_PTP_TSTAMP_OUT;
    output [15:0] TX_PTP_TSTAMP_TAG_OUT;
    output TX_PTP_TSTAMP_VALID_OUT;
    output TX_RDYOUT;
    output [15:0] TX_SERDES_ALT_DATA0;
    output [15:0] TX_SERDES_ALT_DATA1;
    output [15:0] TX_SERDES_ALT_DATA2;
    output [15:0] TX_SERDES_ALT_DATA3;
    output [63:0] TX_SERDES_DATA0;
    output [63:0] TX_SERDES_DATA1;
    output [63:0] TX_SERDES_DATA2;
    output [63:0] TX_SERDES_DATA3;
    output [31:0] TX_SERDES_DATA4;
    output [31:0] TX_SERDES_DATA5;
    output [31:0] TX_SERDES_DATA6;
    output [31:0] TX_SERDES_DATA7;
    output [31:0] TX_SERDES_DATA8;
    output [31:0] TX_SERDES_DATA9;
    output TX_UNFOUT;
    input CTL_CAUI4_MODE;
    input CTL_RSFEC_ENABLE_TRANSCODER_BYPASS_MODE;
    input CTL_RSFEC_IEEE_ERROR_INDICATION_MODE;
    input CTL_RX_CHECK_ETYPE_GCP;
    input CTL_RX_CHECK_ETYPE_GPP;
    input CTL_RX_CHECK_ETYPE_PCP;
    input CTL_RX_CHECK_ETYPE_PPP;
    input CTL_RX_CHECK_MCAST_GCP;
    input CTL_RX_CHECK_MCAST_GPP;
    input CTL_RX_CHECK_MCAST_PCP;
    input CTL_RX_CHECK_MCAST_PPP;
    input CTL_RX_CHECK_OPCODE_GCP;
    input CTL_RX_CHECK_OPCODE_GPP;
    input CTL_RX_CHECK_OPCODE_PCP;
    input CTL_RX_CHECK_OPCODE_PPP;
    input CTL_RX_CHECK_SA_GCP;
    input CTL_RX_CHECK_SA_GPP;
    input CTL_RX_CHECK_SA_PCP;
    input CTL_RX_CHECK_SA_PPP;
    input CTL_RX_CHECK_UCAST_GCP;
    input CTL_RX_CHECK_UCAST_GPP;
    input CTL_RX_CHECK_UCAST_PCP;
    input CTL_RX_CHECK_UCAST_PPP;
    input CTL_RX_ENABLE;
    input CTL_RX_ENABLE_GCP;
    input CTL_RX_ENABLE_GPP;
    input CTL_RX_ENABLE_PCP;
    input CTL_RX_ENABLE_PPP;
    input CTL_RX_FORCE_RESYNC;
    input [8:0] CTL_RX_PAUSE_ACK;
    input [8:0] CTL_RX_PAUSE_ENABLE;
    input CTL_RX_RSFEC_ENABLE;
    input CTL_RX_RSFEC_ENABLE_CORRECTION;
    input CTL_RX_RSFEC_ENABLE_INDICATION;
    input [79:0] CTL_RX_SYSTEMTIMERIN;
    input CTL_RX_TEST_PATTERN;
    input CTL_TX_ENABLE;
    input CTL_TX_LANE0_VLM_BIP7_OVERRIDE;
    input [7:0] CTL_TX_LANE0_VLM_BIP7_OVERRIDE_VALUE;
    input [8:0] CTL_TX_PAUSE_ENABLE;
    input [15:0] CTL_TX_PAUSE_QUANTA0;
    input [15:0] CTL_TX_PAUSE_QUANTA1;
    input [15:0] CTL_TX_PAUSE_QUANTA2;
    input [15:0] CTL_TX_PAUSE_QUANTA3;
    input [15:0] CTL_TX_PAUSE_QUANTA4;
    input [15:0] CTL_TX_PAUSE_QUANTA5;
    input [15:0] CTL_TX_PAUSE_QUANTA6;
    input [15:0] CTL_TX_PAUSE_QUANTA7;
    input [15:0] CTL_TX_PAUSE_QUANTA8;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER0;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER1;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER2;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER3;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER4;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER5;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER6;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER7;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER8;
    input [8:0] CTL_TX_PAUSE_REQ;
    input CTL_TX_PTP_VLANE_ADJUST_MODE;
    input CTL_TX_RESEND_PAUSE;
    input CTL_TX_RSFEC_ENABLE;
    input CTL_TX_SEND_IDLE;
    input CTL_TX_SEND_LFI;
    input CTL_TX_SEND_RFI;
    input [79:0] CTL_TX_SYSTEMTIMERIN;
    input CTL_TX_TEST_PATTERN;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input [329:0] RSFEC_BYPASS_RX_DIN;
    input RSFEC_BYPASS_RX_DIN_CW_START;
    input [329:0] RSFEC_BYPASS_TX_DIN;
    input RSFEC_BYPASS_TX_DIN_CW_START;
    input RX_CLK;
    input RX_RESET;
    input [15:0] RX_SERDES_ALT_DATA0;
    input [15:0] RX_SERDES_ALT_DATA1;
    input [15:0] RX_SERDES_ALT_DATA2;
    input [15:0] RX_SERDES_ALT_DATA3;
    input [9:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA0;
    input [63:0] RX_SERDES_DATA1;
    input [63:0] RX_SERDES_DATA2;
    input [63:0] RX_SERDES_DATA3;
    input [31:0] RX_SERDES_DATA4;
    input [31:0] RX_SERDES_DATA5;
    input [31:0] RX_SERDES_DATA6;
    input [31:0] RX_SERDES_DATA7;
    input [31:0] RX_SERDES_DATA8;
    input [31:0] RX_SERDES_DATA9;
    input [9:0] RX_SERDES_RESET;
    input TX_CLK;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input [55:0] TX_PREIN;
    input [1:0] TX_PTP_1588OP_IN;
    input [15:0] TX_PTP_CHKSUM_OFFSET_IN;
    input [63:0] TX_PTP_RXTSTAMP_IN;
    input [15:0] TX_PTP_TAG_FIELD_IN;
    input [15:0] TX_PTP_TSTAMP_OFFSET_IN;
    input TX_PTP_UPD_CHKSUM_IN;
    input TX_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module GTHE3_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'hF800;
    parameter [15:0] ADAPT_CFG1 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h20F8;
    parameter [15:0] CPLL_CFG1 = 16'hA494;
    parameter [15:0] CPLL_CFG2 = 16'hF001;
    parameter [5:0] CPLL_CFG3 = 6'h00;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [7:0] CPLL_INIT_CFG1 = 8'h00;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DFE_D_X_REL_POS = 1'b0;
    parameter [0:0] DFE_VCM_COMP_EN = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [10:0] EVODD_PHI_CFG = 11'b00000000000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] GM_BIAS_SELECT = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [2:0] PCS_RSVD1 = 3'b000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [1:0] PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [15:0] PMA_RSV1 = 16'h0000;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0000;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG1 = 16'h0080;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h07E6;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG4 = 16'h0000;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG5 = 16'h0000;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h0000;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h5080;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h07E0;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h7C42;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h4000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0060;
    parameter [15:0] RXCFOK_CFG2 = 16'h000E;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0032;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_CFG0 = 16'h0A00;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h7840;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h8000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h8000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_VP_CFG0 = 16'hAA00;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0033;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "Sigcfg_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h8000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0002;
    parameter [8:0] RXOOB_CFG = 9'b000000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h6622;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] RXPI_CFG0 = 2'b00;
    parameter [1:0] RXPI_CFG1 = 2'b00;
    parameter [1:0] RXPI_CFG2 = 2'b00;
    parameter [1:0] RXPI_CFG3 = 2'b00;
    parameter [0:0] RXPI_CFG4 = 1'b0;
    parameter [0:0] RXPI_CFG5 = 1'b1;
    parameter [2:0] RXPI_CFG6 = 3'b000;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h0AD4;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter [7:0] RX_CTLE3_LPF = 8'b00000000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [3:0] RX_DFELPM_CFG0 = 4'b0110;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter [2:0] RX_DFE_AGC_CFG1 = 3'b100;
    parameter [1:0] RX_DFE_KL_LPM_KH_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KH_CFG1 = 3'b010;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_HI_LR = 1'b0;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter real RX_PROGDIV_CFG = 4.0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter [1:0] RX_SUM_RES_CTRL = 2'b00;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b0000;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b000;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [0:0] RX_WIDEMODE_CDR = 1'b0;
    parameter RX_XCLK_SEL = "RXDES";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [0:0] SIM_TX_EIDLE_DRIVE_LEVEL = 1'b0;
    parameter integer SIM_VERSION = 2;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATUR_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter [3:0] TXDRVBIAS_N = 4'b1010;
    parameter [3:0] TXDRVBIAS_P = 4'b1100;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h2020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0001;
    parameter [15:0] TXPH_CFG = 16'h0980;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DCD_CFG = 6'b000010;
    parameter [0:0] TX_DCD_EN = 1'b0;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_EML_PHI_TUNE = 1'b0;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [2:0] TX_MODE_SEL = 3'b000;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 4.0;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [1:0] WB_MODE = 2'b00;
    output [2:0] BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output [2:0] BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [16:0] DMONITOROUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [11:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [7:0] PINRSRVDAS;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output [6:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [8:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input EVODDPHICALDONE;
    input EVODDPHICALSTART;
    input EVODDPHIDRDEN;
    input EVODDPHIDWREN;
    input EVODDPHIXRDEN;
    input EVODDPHIXWREN;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input [2:0] LOOPBACK;
    input LPBKRXTXSEREN;
    input LPBKTXRXSEREN;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input QPLL0CLK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RSTCLKENTX;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input [1:0] RXDFEAGCCTRL;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input [3:0] RXOSINTCFG;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input RXQPIEN;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input [2:0] TXBUFDIFFCTRL;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDEEMPH;
    input TXDETECTRX;
    input [3:0] TXDIFFCTRL;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPRECURSORINV;
    input TXPROGDIVRESET;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTHE3_COMMON (...);
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [9:0] BIAS_CFG_RSVD = 10'b0000000000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0004;
    parameter [15:0] QPLL0_CFG0 = 16'h3018;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0000;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0000;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0009;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h01E8;
    parameter [9:0] QPLL0_LPF = 10'b1111111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter integer QPLL0_REFCLK_DIV = 2;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'b0000000000000000;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] QPLL1_CFG0 = 16'h3018;
    parameter [15:0] QPLL1_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0000;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0000;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0009;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1111111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter integer QPLL1_REFCLK_DIV = 2;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'b0000000000000000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_EN = 1'b1;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0DATA1_0 = 16'b0000000000000000;
    parameter [8:0] SDM0DATA1_1 = 9'b000000000;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [0:0] SDM0_DATA_PIN_SEL = 1'b0;
    parameter [0:0] SDM0_WIDTH_PIN_SEL = 1'b0;
    parameter [15:0] SDM1DATA1_0 = 16'b0000000000000000;
    parameter [8:0] SDM1DATA1_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter [0:0] SDM1_DATA_PIN_SEL = 1'b0;
    parameter [0:0] SDM1_WIDTH_PIN_SEL = 1'b0;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer SIM_VERSION = 2;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0_SEL;
    output [1:0] RXRECCLK1_SEL;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [8:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
endmodule

module GTHE4_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_RXTERMINATION = 1'b1;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter [0:0] CAPBYPASS_FORCE = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter [0:0] CFOK_PWRSVE_EN = 1'b1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h2424;
    parameter [15:0] CKCAL1_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter [15:0] CKCAL_RSVD0 = 16'h4000;
    parameter [15:0] CKCAL_RSVD1 = 16'h0000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h01FA;
    parameter [15:0] CPLL_CFG1 = 16'h24A9;
    parameter [15:0] CPLL_CFG2 = 16'h6807;
    parameter [15:0] CPLL_CFG3 = 16'h0000;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DELAY_ELEC = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h800;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [2:0] LPBK_BIAS_CTRL = 3'b000;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter [2:0] LPBK_IND_CTRL0 = 3'b000;
    parameter [2:0] LPBK_IND_CTRL1 = 3'b000;
    parameter [2:0] LPBK_IND_CTRL2 = 3'b000;
    parameter [3:0] LPBK_RG_CTRL = 4'b0000;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'b00000;
    parameter [5:0] PCIE3_CLK_COR_FULL_THRSH = 6'b010000;
    parameter [4:0] PCIE3_CLK_COR_MAX_LAT = 5'b01000;
    parameter [4:0] PCIE3_CLK_COR_MIN_LAT = 5'b00100;
    parameter [5:0] PCIE3_CLK_COR_THRSH_TIMER = 6'b001000;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN4 = 2'h0;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0;
    parameter [0:0] RCLK_SIPO_INV_EN = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [2:0] RTX_BUF_CML_CTRL = 3'b010;
    parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0003;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0003;
    parameter [15:0] RXCDR_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h0164;
    parameter [9:0] RXCDR_CFG2_GEN2 = 10'h164;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0034;
    parameter [15:0] RXCDR_CFG2_GEN4 = 16'h0034;
    parameter [15:0] RXCDR_CFG3 = 16'h0024;
    parameter [5:0] RXCDR_CFG3_GEN2 = 6'h24;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0024;
    parameter [15:0] RXCDR_CFG3_GEN4 = 16'h0024;
    parameter [15:0] RXCDR_CFG4 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG5 = 16'hB46B;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h146B;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h0000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0002;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_KH_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG3 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0002;
    parameter [0:0] RXDFE_PWR_SAVING = 1'b0;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_UT_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h1000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000110000;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [0:0] RXPI_AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [15:0] RXPI_CFG0 = 16'h0002;
    parameter [15:0] RXPI_CFG1 = 16'b0000000000000000;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [1:0] RXPI_SEL_LC = 2'b00;
    parameter [1:0] RXPI_STARTCODE = 2'b00;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter [0:0] RXREFCLKDIV2_SEL = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h12B0;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 12;
    parameter [7:0] RX_CTLE3_LPF = 8'b00000000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b011;
    parameter integer RX_DFELPM_CFG0 = 0;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b1;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 4;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [0:0] RX_DIV2_MODE_B = 1'b0;
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter [0:0] RX_EN_HI_LR = 1'b1;
    parameter [8:0] RX_EXT_RL_CTRL = 9'b000000000;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] RX_PMA_RSV0 = 16'h0000;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b1001;
    parameter [3:0] RX_SUM_RESLOAD_CTRL = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b1010;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b101;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter [0:0] SAMPLE_CLK_PHASE = 1'b0;
    parameter [0:0] SAS_12G_MODE = 1'b0;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
    parameter [0:0] SRSTMODE = 1'b0;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATURE_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter [3:0] TXDRVBIAS_N = 4'b1010;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h6020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0002;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] TXPI_CFG = 16'h0000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter [0:0] TXPI_PPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXREFCLKDIV2_SEL = 1'b0;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [5:0] TX_DEEMPH2 = 6'b000000;
    parameter [5:0] TX_DEEMPH3 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter integer TX_DRVMUX_CTRL = 2;
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h003F;
    parameter [15:0] TX_PHICAL_CFG2 = 16'h0000;
    parameter integer TX_PI_BIASSET = 0;
    parameter [1:0] TX_PI_IBIAS_MID = 2'b00;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] TX_PMA_RSV0 = 16'h0008;
    parameter integer TX_PREDRV_CTRL = 2;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 3;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter [1:0] TX_SW_MEAS = 2'b00;
    parameter [2:0] TX_VREG_CTRL = 3'b000;
    parameter [0:0] TX_VREG_PDB = 1'b0;
    parameter [1:0] TX_VREG_VREFSEL = 2'b00;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USB_BOTH_BURST_IDLE = 1'b0;
    parameter [6:0] USB_BURSTMAX_U3WAKE = 7'b1111111;
    parameter [6:0] USB_BURSTMIN_U3WAKE = 7'b1100011;
    parameter [0:0] USB_CLK_COR_EQ_EN = 1'b0;
    parameter [0:0] USB_EXT_CNTL = 1'b1;
    parameter [9:0] USB_IDLEMAX_POLLING = 10'b1010111011;
    parameter [9:0] USB_IDLEMIN_POLLING = 10'b0100101011;
    parameter [8:0] USB_LFPSPING_BURST = 9'b000000101;
    parameter [8:0] USB_LFPSPOLLING_BURST = 9'b000110001;
    parameter [8:0] USB_LFPSPOLLING_IDLE_MS = 9'b000000100;
    parameter [8:0] USB_LFPSU1EXIT_BURST = 9'b000011101;
    parameter [8:0] USB_LFPSU2LPEXIT_BURST_MS = 9'b001100011;
    parameter [8:0] USB_LFPSU3WAKE_BURST_MS = 9'b111110011;
    parameter [3:0] USB_LFPS_TPERIOD = 4'b0011;
    parameter [0:0] USB_LFPS_TPERIOD_ACCURATE = 1'b1;
    parameter [0:0] USB_MODE = 1'b0;
    parameter [0:0] USB_PCIE_ERR_REP_DIS = 1'b0;
    parameter integer USB_PING_SATA_MAX_INIT = 21;
    parameter integer USB_PING_SATA_MIN_INIT = 12;
    parameter integer USB_POLL_SATA_MAX_BURST = 8;
    parameter integer USB_POLL_SATA_MIN_BURST = 4;
    parameter [0:0] USB_RAW_ELEC = 1'b0;
    parameter [0:0] USB_RXIDLE_P0_CTRL = 1'b1;
    parameter [0:0] USB_TXIDLE_TUNE_ENABLE = 1'b1;
    parameter integer USB_U1_SATA_MAX_WAKE = 7;
    parameter integer USB_U1_SATA_MIN_WAKE = 4;
    parameter integer USB_U2_SAS_MAX_COM = 64;
    parameter integer USB_U2_SAS_MIN_COM = 36;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [0:0] Y_ALL_MODE = 1'b0;
    output BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [15:0] DMONITOROUT;
    output DMONITOROUTCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [15:0] PINRSRVDAS;
    output POWERPRESENT;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output RXLFPSTRESETDET;
    output RXLFPSU2LPEXITDET;
    output RXLFPSU3WAKEDET;
    output [7:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLFREQLOCK;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input FREQOS;
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTRXRESETSEL;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTTXRESETSEL;
    input INCPCTRL;
    input [2:0] LOOPBACK;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input QPLL0CLK;
    input QPLL0FREQLOCK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1FREQLOCK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXAFECFOKEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input [6:0] RXCKCALSTART;
    input RXCOMMADETEN;
    input [1:0] RXDFEAGCCTRL;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input [3:0] RXDFECFOKFCNUM;
    input RXDFECFOKFEN;
    input RXDFECFOKFPULSE;
    input RXDFECFOKHOLD;
    input RXDFECFOKOVREN;
    input RXDFEKHHOLD;
    input RXDFEKHOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXEQTRAINING;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input RXQPIEN;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXTERMINATION;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input [1:0] TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input TXLFPSTRESET;
    input TXLFPSU2LPEXIT;
    input TXLFPSU3WAKE;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input TXMUXDCDEXHOLD;
    input TXMUXDCDORWREN;
    input TXONESZEROS;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input TXQPIBIASEN;
    input TXQPIWEAKPUP;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTHE4_COMMON (...);
    parameter [0:0] AEN_QPLL0_FBDIV = 1'b1;
    parameter [0:0] AEN_QPLL1_FBDIV = 1'b1;
    parameter [0:0] AEN_SDM0TOGGLE = 1'b0;
    parameter [0:0] AEN_SDM1TOGGLE = 1'b0;
    parameter [0:0] A_SDM0TOGGLE = 1'b0;
    parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000;
    parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000;
    parameter [0:0] A_SDM1TOGGLE = 1'b0;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [15:0] BIAS_CFG_RSVD = 16'h0000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0000;
    parameter [15:0] PPF0_CFG = 16'h0F00;
    parameter [15:0] PPF1_CFG = 16'h0F00;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h391C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0F80;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0002;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1011111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL0_PCI_EN = 1'b0;
    parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL0_REFCLK_DIV = 1;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h691C;
    parameter [15:0] QPLL1_CFG1 = 16'h0020;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0F80;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0002;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1011111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL1_PCI_EN = 1'b0;
    parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL1_REFCLK_DIV = 1;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_ENB = 1'b0;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0SEL;
    output [1:0] RXRECCLK1SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    output [9:0] TCONGPO;
    output TCONRSVDOUT0;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [15:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [2:0] PCIERATEQPLL0;
    input [2:0] PCIERATEQPLL1;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input [7:0] QPLL0FBDIV;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input [7:0] QPLL1FBDIV;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input SDM0TOGGLE;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input SDM1TOGGLE;
    input [1:0] SDM1WIDTH;
    input [9:0] TCONGPI;
    input TCONPOWERUP;
    input [1:0] TCONRESET;
    input [1:0] TCONRSVDIN1;
endmodule

module GTYE3_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'b0000000000000000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter [0:0] CAPBYPASS_FORCE = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h0000;
    parameter [15:0] CKCAL1_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter [15:0] CKCAL_RSVD0 = 16'h0000;
    parameter [15:0] CKCAL_RSVD1 = 16'h0000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h20F8;
    parameter [15:0] CPLL_CFG1 = 16'hA494;
    parameter [15:0] CPLL_CFG2 = 16'hF001;
    parameter [5:0] CPLL_CFG3 = 6'h00;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [7:0] CPLL_INIT_CFG1 = 8'h00;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DFE_D_X_REL_POS = 1'b0;
    parameter [0:0] DFE_VCM_COMP_EN = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter [10:0] EVODD_PHI_CFG = 11'b00000000000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] GM_BIAS_SELECT = 1'b0;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [15:0] LOOP0_CFG = 16'h0000;
    parameter [15:0] LOOP10_CFG = 16'h0000;
    parameter [15:0] LOOP11_CFG = 16'h0000;
    parameter [15:0] LOOP12_CFG = 16'h0000;
    parameter [15:0] LOOP13_CFG = 16'h0000;
    parameter [15:0] LOOP1_CFG = 16'h0000;
    parameter [15:0] LOOP2_CFG = 16'h0000;
    parameter [15:0] LOOP3_CFG = 16'h0000;
    parameter [15:0] LOOP4_CFG = 16'h0000;
    parameter [15:0] LOOP5_CFG = 16'h0000;
    parameter [15:0] LOOP6_CFG = 16'h0000;
    parameter [15:0] LOOP7_CFG = 16'h0000;
    parameter [15:0] LOOP8_CFG = 16'h0000;
    parameter [15:0] LOOP9_CFG = 16'h0000;
    parameter [2:0] LPBK_BIAS_CTRL = 3'b000;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter [3:0] LPBK_RG_CTRL = 4'b0000;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [2:0] PCS_RSVD1 = 3'b000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [1:0] PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [15:0] PMA_RSV0 = 16'h0000;
    parameter [15:0] PMA_RSV1 = 16'h0000;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0000;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG1 = 16'h0300;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0300;
    parameter [15:0] RXCDR_CFG2 = 16'h0060;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0060;
    parameter [15:0] RXCDR_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG4 = 16'h0002;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h0002;
    parameter [15:0] RXCDR_CFG5 = 16'h0000;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h0000;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0001;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [1:0] RXCFOKDONE_SRC = 2'b00;
    parameter [15:0] RXCFOK_CFG0 = 16'h3E00;
    parameter [15:0] RXCFOK_CFG1 = 16'h0042;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4C00;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h1E00;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h1900;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0200;
    parameter [0:0] RXDFE_PWR_SAVING = 1'b0;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h0200;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0400;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [0:0] RXPI_AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [15:0] RXPI_CFG = 16'h0100;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [15:0] RXPI_RSV0 = 16'h0000;
    parameter [1:0] RXPI_SEL_LC = 2'b00;
    parameter [1:0] RXPI_STARTCODE = 2'b00;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h1534;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 10;
    parameter [0:0] RX_CTLE1_KHKL = 1'b0;
    parameter [0:0] RX_CTLE2_KHKL = 1'b0;
    parameter [0:0] RX_CTLE3_AGC = 1'b0;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b010;
    parameter integer RX_DFELPM_CFG0 = 6;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 2;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [0:0] RX_DIV2_MODE_B = 1'b0;
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter [0:0] RX_EN_HI_LR = 1'b0;
    parameter [8:0] RX_EXT_RL_CTRL = 9'b000000000;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b1000;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b101;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [0:0] SIM_TX_EIDLE_DRIVE_LEVEL = 1'b0;
    parameter integer SIM_VERSION = 2;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATURE_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h2020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0001;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [15:0] TXPI_RSV0 = 16'h0000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter [0:0] TX_CLKREG_PDB = 1'b0;
    parameter [2:0] TX_CLKREG_SET = 3'b000;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DCD_CFG = 6'b000010;
    parameter [0:0] TX_DCD_EN = 1'b0;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter integer TX_DRVMUX_CTRL = 2;
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_EML_PHI_TUNE = 1'b0;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [2:0] TX_MODE_SEL = 3'b000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h7E00;
    parameter [15:0] TX_PHICAL_CFG2 = 16'h0000;
    parameter integer TX_PI_BIASSET = 0;
    parameter [15:0] TX_PI_CFG0 = 16'h0000;
    parameter [15:0] TX_PI_CFG1 = 16'h0000;
    parameter [0:0] TX_PI_DIV2_MODE_B = 1'b0;
    parameter [0:0] TX_PI_SEL_QPLL0 = 1'b0;
    parameter [0:0] TX_PI_SEL_QPLL1 = 1'b0;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter integer TX_PREDRV_CTRL = 2;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 4;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output [2:0] BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output [2:0] BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [16:0] DMONITOROUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output GTYTXN;
    output GTYTXP;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [7:0] PINRSRVDAS;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output [6:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input ELPCALDVORWREN;
    input ELPCALPAORWREN;
    input EVODDPHICALDONE;
    input EVODDPHICALSTART;
    input EVODDPHIDRDEN;
    input EVODDPHIDWREN;
    input EVODDPHIXRDEN;
    input EVODDPHIXWREN;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTYRXN;
    input GTYRXP;
    input [2:0] LOOPBACK;
    input [15:0] LOOPRSVD;
    input LPBKRXTXSEREN;
    input LPBKTXRXSEREN;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input QPLL0CLK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RSTCLKENTX;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input RXCOMMADETEN;
    input RXDCCFORCESTART;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input [3:0] RXOSINTCFG;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input [2:0] TXBUFDIFFCTRL;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXELFORCESTART;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTYE3_COMMON (...);
    parameter [15:0] A_SDM1DATA1_0 = 16'b0000000000000000;
    parameter [8:0] A_SDM1DATA1_1 = 9'b000000000;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [9:0] BIAS_CFG_RSVD = 10'b0000000000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0004;
    parameter [15:0] PPF0_CFG = 16'h0FFF;
    parameter [15:0] PPF1_CFG = 16'h0FFF;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h301C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0780;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0780;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0021;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1111111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter integer QPLL0_REFCLK_DIV = 2;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h301C;
    parameter [15:0] QPLL1_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0780;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0780;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0021;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1111111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter integer QPLL1_REFCLK_DIV = 2;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_EN = 1'b1;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer SIM_VERSION = 2;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0_SEL;
    output [1:0] RXRECCLK1_SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input [1:0] SDM1WIDTH;
endmodule

module GTYE4_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_RXTERMINATION = 1'b1;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter [0:0] CFOK_PWRSVE_EN = 1'b1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h2424;
    parameter [15:0] CKCAL1_CFG_0 = 16'b1100000011000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0101000011000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b1100000011000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b1000000011000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h01FA;
    parameter [15:0] CPLL_CFG1 = 16'h24A9;
    parameter [15:0] CPLL_CFG2 = 16'h6807;
    parameter [15:0] CPLL_CFG3 = 16'h0000;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DELAY_ELEC = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h800;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter integer EYESCAN_VP_RANGE = 0;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter integer LPBK_BIAS_CTRL = 4;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter integer LPBK_IND_CTRL0 = 5;
    parameter integer LPBK_IND_CTRL1 = 5;
    parameter integer LPBK_IND_CTRL2 = 5;
    parameter integer LPBK_RG_CTRL = 2;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'b00000;
    parameter [5:0] PCIE3_CLK_COR_FULL_THRSH = 6'b010000;
    parameter [4:0] PCIE3_CLK_COR_MAX_LAT = 5'b01000;
    parameter [4:0] PCIE3_CLK_COR_MIN_LAT = 5'b00100;
    parameter [5:0] PCIE3_CLK_COR_THRSH_TIMER = 6'b001000;
    parameter PCIE_64B_DYN_CLKSW_DIS = "FALSE";
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter PCIE_GEN4_64BIT_INT_EN = "FALSE";
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN4 = 2'h0;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'h0000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0;
    parameter [0:0] RCLK_SIPO_INV_EN = 1'b0;
    parameter [2:0] RTX_BUF_CML_CTRL = 3'b010;
    parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b10000;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0003;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0003;
    parameter [15:0] RXCDR_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h0164;
    parameter [9:0] RXCDR_CFG2_GEN2 = 10'h164;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0034;
    parameter [15:0] RXCDR_CFG2_GEN4 = 16'h0034;
    parameter [15:0] RXCDR_CFG3 = 16'h0024;
    parameter [5:0] RXCDR_CFG3_GEN2 = 6'h24;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0024;
    parameter [15:0] RXCDR_CFG3_GEN4 = 16'h0024;
    parameter [15:0] RXCDR_CFG4 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG5 = 16'hB46B;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h146B;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h0000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0002;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_KH_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG3 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_UT_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h1000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000110000;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] RXPI_CFG0 = 16'h0102;
    parameter [15:0] RXPI_CFG1 = 16'b0000000001010100;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter [0:0] RXREFCLKDIV2_SEL = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h12B0;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 12;
    parameter [0:0] RX_CTLE_PWR_SAVING = 1'b0;
    parameter [3:0] RX_CTLE_RES_CTRL = 4'b0000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b100;
    parameter integer RX_DFELPM_CFG0 = 0;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b1;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 4;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter integer RX_EN_SUM_RCAL_B = 0;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b10;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] RX_I2V_FILTER_EN = 1'b1;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] RX_PMA_RSV0 = 16'h000F;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter integer RX_SUM_DEGEN_AVTT_OVERITE = 0;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter integer RX_SUM_PWR_SAVING = 0;
    parameter [3:0] RX_SUM_RES_CTRL = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b0011;
    parameter [0:0] RX_SUM_VCM_BIAS_TUNE_EN = 1'b1;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b010;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter [0:0] SAMPLE_CLK_PHASE = 1'b0;
    parameter [0:0] SAS_12G_MODE = 1'b0;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [0:0] SRSTMODE = 1'b0;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter integer TXDRV_FREQBAND = 0;
    parameter [15:0] TXFE_CFG0 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG1 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG2 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG3 = 16'b0000000000000000;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h6020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0002;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] TXPI_CFG0 = 16'b0000000100000000;
    parameter [15:0] TXPI_CFG1 = 16'b0000000000000000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_PPM = 1'b0;
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXREFCLKDIV2_SEL = 1'b0;
    parameter integer TXSWBST_BST = 1;
    parameter integer TXSWBST_EN = 0;
    parameter integer TXSWBST_MAG = 6;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [5:0] TX_DEEMPH2 = 6'b000000;
    parameter [5:0] TX_DEEMPH3 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h003F;
    parameter integer TX_PI_BIASSET = 0;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] TX_PMA_RSV0 = 16'h0000;
    parameter [15:0] TX_PMA_RSV1 = 16'h0000;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 3;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [1:0] TX_SW_MEAS = 2'b00;
    parameter [2:0] TX_VREG_CTRL = 3'b000;
    parameter [0:0] TX_VREG_PDB = 1'b0;
    parameter [1:0] TX_VREG_VREFSEL = 2'b00;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USB_BOTH_BURST_IDLE = 1'b0;
    parameter [6:0] USB_BURSTMAX_U3WAKE = 7'b1111111;
    parameter [6:0] USB_BURSTMIN_U3WAKE = 7'b1100011;
    parameter [0:0] USB_CLK_COR_EQ_EN = 1'b0;
    parameter [0:0] USB_EXT_CNTL = 1'b1;
    parameter [9:0] USB_IDLEMAX_POLLING = 10'b1010111011;
    parameter [9:0] USB_IDLEMIN_POLLING = 10'b0100101011;
    parameter [8:0] USB_LFPSPING_BURST = 9'b000000101;
    parameter [8:0] USB_LFPSPOLLING_BURST = 9'b000110001;
    parameter [8:0] USB_LFPSPOLLING_IDLE_MS = 9'b000000100;
    parameter [8:0] USB_LFPSU1EXIT_BURST = 9'b000011101;
    parameter [8:0] USB_LFPSU2LPEXIT_BURST_MS = 9'b001100011;
    parameter [8:0] USB_LFPSU3WAKE_BURST_MS = 9'b111110011;
    parameter [3:0] USB_LFPS_TPERIOD = 4'b0011;
    parameter [0:0] USB_LFPS_TPERIOD_ACCURATE = 1'b1;
    parameter [0:0] USB_MODE = 1'b0;
    parameter [0:0] USB_PCIE_ERR_REP_DIS = 1'b0;
    parameter integer USB_PING_SATA_MAX_INIT = 21;
    parameter integer USB_PING_SATA_MIN_INIT = 12;
    parameter integer USB_POLL_SATA_MAX_BURST = 8;
    parameter integer USB_POLL_SATA_MIN_BURST = 4;
    parameter [0:0] USB_RAW_ELEC = 1'b0;
    parameter [0:0] USB_RXIDLE_P0_CTRL = 1'b1;
    parameter [0:0] USB_TXIDLE_TUNE_ENABLE = 1'b1;
    parameter integer USB_U1_SATA_MAX_WAKE = 7;
    parameter integer USB_U1_SATA_MIN_WAKE = 4;
    parameter integer USB_U2_SAS_MAX_COM = 64;
    parameter integer USB_U2_SAS_MIN_COM = 36;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [0:0] Y_ALL_MODE = 1'b0;
    output BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [15:0] DMONITOROUT;
    output DMONITOROUTCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output GTYTXN;
    output GTYTXP;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [15:0] PINRSRVDAS;
    output POWERPRESENT;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output RXLFPSTRESETDET;
    output RXLFPSU2LPEXITDET;
    output RXLFPSU3WAKEDET;
    output [7:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLFREQLOCK;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input FREQOS;
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTRXRESETSEL;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTTXRESETSEL;
    input GTYRXN;
    input GTYRXP;
    input INCPCTRL;
    input [2:0] LOOPBACK;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input QPLL0CLK;
    input QPLL0FREQLOCK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1FREQLOCK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXAFECFOKEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input [6:0] RXCKCALSTART;
    input RXCOMMADETEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input [3:0] RXDFECFOKFCNUM;
    input RXDFECFOKFEN;
    input RXDFECFOKFPULSE;
    input RXDFECFOKHOLD;
    input RXDFECFOKOVREN;
    input RXDFEKHHOLD;
    input RXDFEKHOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXEQTRAINING;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXTERMINATION;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input [1:0] TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input TXLFPSTRESET;
    input TXLFPSU2LPEXIT;
    input TXLFPSU3WAKE;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input TXMUXDCDEXHOLD;
    input TXMUXDCDORWREN;
    input TXONESZEROS;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTYE4_COMMON (...);
    parameter [0:0] AEN_QPLL0_FBDIV = 1'b1;
    parameter [0:0] AEN_QPLL1_FBDIV = 1'b1;
    parameter [0:0] AEN_SDM0TOGGLE = 1'b0;
    parameter [0:0] AEN_SDM1TOGGLE = 1'b0;
    parameter [0:0] A_SDM0TOGGLE = 1'b0;
    parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000;
    parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000;
    parameter [0:0] A_SDM1TOGGLE = 1'b0;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [15:0] BIAS_CFG_RSVD = 16'h0000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0000;
    parameter [15:0] PPF0_CFG = 16'h0F00;
    parameter [15:0] PPF1_CFG = 16'h0F00;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h391C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0F80;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0002;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1011111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL0_PCI_EN = 1'b0;
    parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL0_REFCLK_DIV = 1;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h691C;
    parameter [15:0] QPLL1_CFG1 = 16'h0020;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0F80;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0002;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1011111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL1_PCI_EN = 1'b0;
    parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL1_REFCLK_DIV = 1;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_ENB = 1'b0;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [15:0] UB_CFG0 = 16'h0000;
    parameter [15:0] UB_CFG1 = 16'h0000;
    parameter [15:0] UB_CFG2 = 16'h0000;
    parameter [15:0] UB_CFG3 = 16'h0000;
    parameter [15:0] UB_CFG4 = 16'h0000;
    parameter [15:0] UB_CFG5 = 16'h0400;
    parameter [15:0] UB_CFG6 = 16'h0000;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0SEL;
    output [1:0] RXRECCLK1SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    output [15:0] UBDADDR;
    output UBDEN;
    output [15:0] UBDI;
    output UBDWE;
    output UBMDMTDO;
    output UBRSVDOUT;
    output UBTXUART;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [15:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [2:0] PCIERATEQPLL0;
    input [2:0] PCIERATEQPLL1;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input [7:0] QPLL0FBDIV;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input [7:0] QPLL1FBDIV;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input SDM0TOGGLE;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input SDM1TOGGLE;
    input [1:0] SDM1WIDTH;
    input UBCFGSTREAMEN;
    input [15:0] UBDO;
    input UBDRDY;
    input UBENABLE;
    input [1:0] UBGPI;
    input [1:0] UBINTR;
    input UBIOLMBRST;
    input UBMBRST;
    input UBMDMCAPTURE;
    input UBMDMDBGRST;
    input UBMDMDBGUPDATE;
    input [3:0] UBMDMREGEN;
    input UBMDMSHIFT;
    input UBMDMSYSRST;
    input UBMDMTCK;
    input UBMDMTDI;
endmodule

module IBUFDS_GTE3 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [1:0] REFCLK_HROW_CK_SEL = 2'b00;
    parameter [1:0] REFCLK_ICNTL_RX = 2'b00;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_GTE4 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [1:0] REFCLK_HROW_CK_SEL = 2'b00;
    parameter [1:0] REFCLK_ICNTL_RX = 2'b00;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module ILKN (...);
    parameter BYPASS = "FALSE";
    parameter [1:0] CTL_RX_BURSTMAX = 2'h3;
    parameter [1:0] CTL_RX_CHAN_EXT = 2'h0;
    parameter [3:0] CTL_RX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_RX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter CTL_RX_PACKET_MODE = "TRUE";
    parameter [2:0] CTL_RX_RETRANS_MULT = 3'h0;
    parameter [3:0] CTL_RX_RETRANS_RETRY = 4'h2;
    parameter [15:0] CTL_RX_RETRANS_TIMER1 = 16'h0000;
    parameter [15:0] CTL_RX_RETRANS_TIMER2 = 16'h0008;
    parameter [11:0] CTL_RX_RETRANS_WDOG = 12'h000;
    parameter [7:0] CTL_RX_RETRANS_WRAP_TIMER = 8'h00;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [1:0] CTL_TX_BURSTMAX = 2'h3;
    parameter [2:0] CTL_TX_BURSTSHORT = 3'h1;
    parameter [1:0] CTL_TX_CHAN_EXT = 2'h0;
    parameter CTL_TX_DISABLE_SKIPWORD = "TRUE";
    parameter [6:0] CTL_TX_FC_CALLEN = 7'h00;
    parameter [3:0] CTL_TX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_TX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter [13:0] CTL_TX_RETRANS_DEPTH = 14'h0800;
    parameter [2:0] CTL_TX_RETRANS_MULT = 3'h0;
    parameter [1:0] CTL_TX_RETRANS_RAM_BANKS = 2'h3;
    parameter MODE = "TRUE";
    parameter SIM_VERSION = "2.0";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [65:0] RX_BYPASS_DATAOUT00;
    output [65:0] RX_BYPASS_DATAOUT01;
    output [65:0] RX_BYPASS_DATAOUT02;
    output [65:0] RX_BYPASS_DATAOUT03;
    output [65:0] RX_BYPASS_DATAOUT04;
    output [65:0] RX_BYPASS_DATAOUT05;
    output [65:0] RX_BYPASS_DATAOUT06;
    output [65:0] RX_BYPASS_DATAOUT07;
    output [65:0] RX_BYPASS_DATAOUT08;
    output [65:0] RX_BYPASS_DATAOUT09;
    output [65:0] RX_BYPASS_DATAOUT10;
    output [65:0] RX_BYPASS_DATAOUT11;
    output [11:0] RX_BYPASS_ENAOUT;
    output [11:0] RX_BYPASS_IS_AVAILOUT;
    output [11:0] RX_BYPASS_IS_BADLYFRAMEDOUT;
    output [11:0] RX_BYPASS_IS_OVERFLOWOUT;
    output [11:0] RX_BYPASS_IS_SYNCEDOUT;
    output [11:0] RX_BYPASS_IS_SYNCWORDOUT;
    output [10:0] RX_CHANOUT0;
    output [10:0] RX_CHANOUT1;
    output [10:0] RX_CHANOUT2;
    output [10:0] RX_CHANOUT3;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output RX_OVFOUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [11:0] STAT_RX_BAD_TYPE_ERR;
    output STAT_RX_BURSTMAX_ERR;
    output STAT_RX_BURST_ERR;
    output STAT_RX_CRC24_ERR;
    output [11:0] STAT_RX_CRC32_ERR;
    output [11:0] STAT_RX_CRC32_VALID;
    output [11:0] STAT_RX_DESCRAM_ERR;
    output [11:0] STAT_RX_DIAGWORD_INTFSTAT;
    output [11:0] STAT_RX_DIAGWORD_LANESTAT;
    output [255:0] STAT_RX_FC_STAT;
    output [11:0] STAT_RX_FRAMING_ERR;
    output STAT_RX_MEOP_ERR;
    output [11:0] STAT_RX_MF_ERR;
    output [11:0] STAT_RX_MF_LEN_ERR;
    output [11:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MSOP_ERR;
    output [7:0] STAT_RX_MUBITS;
    output STAT_RX_MUBITS_UPDATED;
    output STAT_RX_OVERFLOW_ERR;
    output STAT_RX_RETRANS_CRC24_ERR;
    output STAT_RX_RETRANS_DISC;
    output [15:0] STAT_RX_RETRANS_LATENCY;
    output STAT_RX_RETRANS_REQ;
    output STAT_RX_RETRANS_RETRY_ERR;
    output [7:0] STAT_RX_RETRANS_SEQ;
    output STAT_RX_RETRANS_SEQ_UPDATED;
    output [2:0] STAT_RX_RETRANS_STATE;
    output [4:0] STAT_RX_RETRANS_SUBSEQ;
    output STAT_RX_RETRANS_WDOG_ERR;
    output STAT_RX_RETRANS_WRAP_ERR;
    output [11:0] STAT_RX_SYNCED;
    output [11:0] STAT_RX_SYNCED_ERR;
    output [11:0] STAT_RX_WORD_SYNC;
    output STAT_TX_BURST_ERR;
    output STAT_TX_ERRINJ_BITERR_DONE;
    output STAT_TX_OVERFLOW_ERR;
    output STAT_TX_RETRANS_BURST_ERR;
    output STAT_TX_RETRANS_BUSY;
    output STAT_TX_RETRANS_RAM_PERROUT;
    output [8:0] STAT_TX_RETRANS_RAM_RADDR;
    output STAT_TX_RETRANS_RAM_RD_B0;
    output STAT_TX_RETRANS_RAM_RD_B1;
    output STAT_TX_RETRANS_RAM_RD_B2;
    output STAT_TX_RETRANS_RAM_RD_B3;
    output [1:0] STAT_TX_RETRANS_RAM_RSEL;
    output [8:0] STAT_TX_RETRANS_RAM_WADDR;
    output [643:0] STAT_TX_RETRANS_RAM_WDATA;
    output STAT_TX_RETRANS_RAM_WE_B0;
    output STAT_TX_RETRANS_RAM_WE_B1;
    output STAT_TX_RETRANS_RAM_WE_B2;
    output STAT_TX_RETRANS_RAM_WE_B3;
    output STAT_TX_UNDERFLOW_ERR;
    output TX_OVFOUT;
    output TX_RDYOUT;
    output [63:0] TX_SERDES_DATA00;
    output [63:0] TX_SERDES_DATA01;
    output [63:0] TX_SERDES_DATA02;
    output [63:0] TX_SERDES_DATA03;
    output [63:0] TX_SERDES_DATA04;
    output [63:0] TX_SERDES_DATA05;
    output [63:0] TX_SERDES_DATA06;
    output [63:0] TX_SERDES_DATA07;
    output [63:0] TX_SERDES_DATA08;
    output [63:0] TX_SERDES_DATA09;
    output [63:0] TX_SERDES_DATA10;
    output [63:0] TX_SERDES_DATA11;
    input CORE_CLK;
    input CTL_RX_FORCE_RESYNC;
    input CTL_RX_RETRANS_ACK;
    input CTL_RX_RETRANS_ENABLE;
    input CTL_RX_RETRANS_ERRIN;
    input CTL_RX_RETRANS_FORCE_REQ;
    input CTL_RX_RETRANS_RESET;
    input CTL_RX_RETRANS_RESET_MODE;
    input CTL_TX_DIAGWORD_INTFSTAT;
    input [11:0] CTL_TX_DIAGWORD_LANESTAT;
    input CTL_TX_ENABLE;
    input CTL_TX_ERRINJ_BITERR_GO;
    input [3:0] CTL_TX_ERRINJ_BITERR_LANE;
    input [255:0] CTL_TX_FC_STAT;
    input [7:0] CTL_TX_MUBITS;
    input CTL_TX_RETRANS_ENABLE;
    input CTL_TX_RETRANS_RAM_PERRIN;
    input [643:0] CTL_TX_RETRANS_RAM_RDATA;
    input CTL_TX_RETRANS_REQ;
    input CTL_TX_RETRANS_REQ_VALID;
    input [11:0] CTL_TX_RLIM_DELTA;
    input CTL_TX_RLIM_ENABLE;
    input [7:0] CTL_TX_RLIM_INTV;
    input [11:0] CTL_TX_RLIM_MAX;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input LBUS_CLK;
    input RX_BYPASS_FORCE_REALIGNIN;
    input RX_BYPASS_RDIN;
    input RX_RESET;
    input [11:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA00;
    input [63:0] RX_SERDES_DATA01;
    input [63:0] RX_SERDES_DATA02;
    input [63:0] RX_SERDES_DATA03;
    input [63:0] RX_SERDES_DATA04;
    input [63:0] RX_SERDES_DATA05;
    input [63:0] RX_SERDES_DATA06;
    input [63:0] RX_SERDES_DATA07;
    input [63:0] RX_SERDES_DATA08;
    input [63:0] RX_SERDES_DATA09;
    input [63:0] RX_SERDES_DATA10;
    input [63:0] RX_SERDES_DATA11;
    input [11:0] RX_SERDES_RESET;
    input TX_BCTLIN0;
    input TX_BCTLIN1;
    input TX_BCTLIN2;
    input TX_BCTLIN3;
    input [11:0] TX_BYPASS_CTRLIN;
    input [63:0] TX_BYPASS_DATAIN00;
    input [63:0] TX_BYPASS_DATAIN01;
    input [63:0] TX_BYPASS_DATAIN02;
    input [63:0] TX_BYPASS_DATAIN03;
    input [63:0] TX_BYPASS_DATAIN04;
    input [63:0] TX_BYPASS_DATAIN05;
    input [63:0] TX_BYPASS_DATAIN06;
    input [63:0] TX_BYPASS_DATAIN07;
    input [63:0] TX_BYPASS_DATAIN08;
    input [63:0] TX_BYPASS_DATAIN09;
    input [63:0] TX_BYPASS_DATAIN10;
    input [63:0] TX_BYPASS_DATAIN11;
    input TX_BYPASS_ENAIN;
    input [7:0] TX_BYPASS_GEARBOX_SEQIN;
    input [3:0] TX_BYPASS_MFRAMER_STATEIN;
    input [10:0] TX_CHANIN0;
    input [10:0] TX_CHANIN1;
    input [10:0] TX_CHANIN2;
    input [10:0] TX_CHANIN3;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input TX_RESET;
    input TX_SERDES_REFCLK;
    input TX_SERDES_REFCLK_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module ILKNE4 (...);
    parameter BYPASS = "FALSE";
    parameter [1:0] CTL_RX_BURSTMAX = 2'h3;
    parameter [1:0] CTL_RX_CHAN_EXT = 2'h0;
    parameter [3:0] CTL_RX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_RX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter CTL_RX_PACKET_MODE = "FALSE";
    parameter [2:0] CTL_RX_RETRANS_MULT = 3'h0;
    parameter [3:0] CTL_RX_RETRANS_RETRY = 4'h2;
    parameter [15:0] CTL_RX_RETRANS_TIMER1 = 16'h0009;
    parameter [15:0] CTL_RX_RETRANS_TIMER2 = 16'h0000;
    parameter [11:0] CTL_RX_RETRANS_WDOG = 12'h000;
    parameter [7:0] CTL_RX_RETRANS_WRAP_TIMER = 8'h00;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [1:0] CTL_TX_BURSTMAX = 2'h3;
    parameter [2:0] CTL_TX_BURSTSHORT = 3'h1;
    parameter [1:0] CTL_TX_CHAN_EXT = 2'h0;
    parameter CTL_TX_DISABLE_SKIPWORD = "FALSE";
    parameter [3:0] CTL_TX_FC_CALLEN = 4'hF;
    parameter [3:0] CTL_TX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_TX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter [13:0] CTL_TX_RETRANS_DEPTH = 14'h0800;
    parameter [2:0] CTL_TX_RETRANS_MULT = 3'h0;
    parameter [1:0] CTL_TX_RETRANS_RAM_BANKS = 2'h3;
    parameter MODE = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [65:0] RX_BYPASS_DATAOUT00;
    output [65:0] RX_BYPASS_DATAOUT01;
    output [65:0] RX_BYPASS_DATAOUT02;
    output [65:0] RX_BYPASS_DATAOUT03;
    output [65:0] RX_BYPASS_DATAOUT04;
    output [65:0] RX_BYPASS_DATAOUT05;
    output [65:0] RX_BYPASS_DATAOUT06;
    output [65:0] RX_BYPASS_DATAOUT07;
    output [65:0] RX_BYPASS_DATAOUT08;
    output [65:0] RX_BYPASS_DATAOUT09;
    output [65:0] RX_BYPASS_DATAOUT10;
    output [65:0] RX_BYPASS_DATAOUT11;
    output [11:0] RX_BYPASS_ENAOUT;
    output [11:0] RX_BYPASS_IS_AVAILOUT;
    output [11:0] RX_BYPASS_IS_BADLYFRAMEDOUT;
    output [11:0] RX_BYPASS_IS_OVERFLOWOUT;
    output [11:0] RX_BYPASS_IS_SYNCEDOUT;
    output [11:0] RX_BYPASS_IS_SYNCWORDOUT;
    output [10:0] RX_CHANOUT0;
    output [10:0] RX_CHANOUT1;
    output [10:0] RX_CHANOUT2;
    output [10:0] RX_CHANOUT3;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output RX_OVFOUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [11:0] STAT_RX_BAD_TYPE_ERR;
    output STAT_RX_BURSTMAX_ERR;
    output STAT_RX_BURST_ERR;
    output STAT_RX_CRC24_ERR;
    output [11:0] STAT_RX_CRC32_ERR;
    output [11:0] STAT_RX_CRC32_VALID;
    output [11:0] STAT_RX_DESCRAM_ERR;
    output [11:0] STAT_RX_DIAGWORD_INTFSTAT;
    output [11:0] STAT_RX_DIAGWORD_LANESTAT;
    output [255:0] STAT_RX_FC_STAT;
    output [11:0] STAT_RX_FRAMING_ERR;
    output STAT_RX_MEOP_ERR;
    output [11:0] STAT_RX_MF_ERR;
    output [11:0] STAT_RX_MF_LEN_ERR;
    output [11:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MSOP_ERR;
    output [7:0] STAT_RX_MUBITS;
    output STAT_RX_MUBITS_UPDATED;
    output STAT_RX_OVERFLOW_ERR;
    output STAT_RX_RETRANS_CRC24_ERR;
    output STAT_RX_RETRANS_DISC;
    output [15:0] STAT_RX_RETRANS_LATENCY;
    output STAT_RX_RETRANS_REQ;
    output STAT_RX_RETRANS_RETRY_ERR;
    output [7:0] STAT_RX_RETRANS_SEQ;
    output STAT_RX_RETRANS_SEQ_UPDATED;
    output [2:0] STAT_RX_RETRANS_STATE;
    output [4:0] STAT_RX_RETRANS_SUBSEQ;
    output STAT_RX_RETRANS_WDOG_ERR;
    output STAT_RX_RETRANS_WRAP_ERR;
    output [11:0] STAT_RX_SYNCED;
    output [11:0] STAT_RX_SYNCED_ERR;
    output [11:0] STAT_RX_WORD_SYNC;
    output STAT_TX_BURST_ERR;
    output STAT_TX_ERRINJ_BITERR_DONE;
    output STAT_TX_OVERFLOW_ERR;
    output STAT_TX_RETRANS_BURST_ERR;
    output STAT_TX_RETRANS_BUSY;
    output STAT_TX_RETRANS_RAM_PERROUT;
    output [8:0] STAT_TX_RETRANS_RAM_RADDR;
    output STAT_TX_RETRANS_RAM_RD_B0;
    output STAT_TX_RETRANS_RAM_RD_B1;
    output STAT_TX_RETRANS_RAM_RD_B2;
    output STAT_TX_RETRANS_RAM_RD_B3;
    output [1:0] STAT_TX_RETRANS_RAM_RSEL;
    output [8:0] STAT_TX_RETRANS_RAM_WADDR;
    output [643:0] STAT_TX_RETRANS_RAM_WDATA;
    output STAT_TX_RETRANS_RAM_WE_B0;
    output STAT_TX_RETRANS_RAM_WE_B1;
    output STAT_TX_RETRANS_RAM_WE_B2;
    output STAT_TX_RETRANS_RAM_WE_B3;
    output STAT_TX_UNDERFLOW_ERR;
    output TX_OVFOUT;
    output TX_RDYOUT;
    output [63:0] TX_SERDES_DATA00;
    output [63:0] TX_SERDES_DATA01;
    output [63:0] TX_SERDES_DATA02;
    output [63:0] TX_SERDES_DATA03;
    output [63:0] TX_SERDES_DATA04;
    output [63:0] TX_SERDES_DATA05;
    output [63:0] TX_SERDES_DATA06;
    output [63:0] TX_SERDES_DATA07;
    output [63:0] TX_SERDES_DATA08;
    output [63:0] TX_SERDES_DATA09;
    output [63:0] TX_SERDES_DATA10;
    output [63:0] TX_SERDES_DATA11;
    input CORE_CLK;
    input CTL_RX_FORCE_RESYNC;
    input CTL_RX_RETRANS_ACK;
    input CTL_RX_RETRANS_ENABLE;
    input CTL_RX_RETRANS_ERRIN;
    input CTL_RX_RETRANS_FORCE_REQ;
    input CTL_RX_RETRANS_RESET;
    input CTL_RX_RETRANS_RESET_MODE;
    input CTL_TX_DIAGWORD_INTFSTAT;
    input [11:0] CTL_TX_DIAGWORD_LANESTAT;
    input CTL_TX_ENABLE;
    input CTL_TX_ERRINJ_BITERR_GO;
    input [3:0] CTL_TX_ERRINJ_BITERR_LANE;
    input [255:0] CTL_TX_FC_STAT;
    input [7:0] CTL_TX_MUBITS;
    input CTL_TX_RETRANS_ENABLE;
    input CTL_TX_RETRANS_RAM_PERRIN;
    input [643:0] CTL_TX_RETRANS_RAM_RDATA;
    input CTL_TX_RETRANS_REQ;
    input CTL_TX_RETRANS_REQ_VALID;
    input [11:0] CTL_TX_RLIM_DELTA;
    input CTL_TX_RLIM_ENABLE;
    input [7:0] CTL_TX_RLIM_INTV;
    input [11:0] CTL_TX_RLIM_MAX;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input LBUS_CLK;
    input RX_BYPASS_FORCE_REALIGNIN;
    input RX_BYPASS_RDIN;
    input RX_RESET;
    input [11:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA00;
    input [63:0] RX_SERDES_DATA01;
    input [63:0] RX_SERDES_DATA02;
    input [63:0] RX_SERDES_DATA03;
    input [63:0] RX_SERDES_DATA04;
    input [63:0] RX_SERDES_DATA05;
    input [63:0] RX_SERDES_DATA06;
    input [63:0] RX_SERDES_DATA07;
    input [63:0] RX_SERDES_DATA08;
    input [63:0] RX_SERDES_DATA09;
    input [63:0] RX_SERDES_DATA10;
    input [63:0] RX_SERDES_DATA11;
    input [11:0] RX_SERDES_RESET;
    input TX_BCTLIN0;
    input TX_BCTLIN1;
    input TX_BCTLIN2;
    input TX_BCTLIN3;
    input [11:0] TX_BYPASS_CTRLIN;
    input [63:0] TX_BYPASS_DATAIN00;
    input [63:0] TX_BYPASS_DATAIN01;
    input [63:0] TX_BYPASS_DATAIN02;
    input [63:0] TX_BYPASS_DATAIN03;
    input [63:0] TX_BYPASS_DATAIN04;
    input [63:0] TX_BYPASS_DATAIN05;
    input [63:0] TX_BYPASS_DATAIN06;
    input [63:0] TX_BYPASS_DATAIN07;
    input [63:0] TX_BYPASS_DATAIN08;
    input [63:0] TX_BYPASS_DATAIN09;
    input [63:0] TX_BYPASS_DATAIN10;
    input [63:0] TX_BYPASS_DATAIN11;
    input TX_BYPASS_ENAIN;
    input [7:0] TX_BYPASS_GEARBOX_SEQIN;
    input [3:0] TX_BYPASS_MFRAMER_STATEIN;
    input [10:0] TX_CHANIN0;
    input [10:0] TX_CHANIN1;
    input [10:0] TX_CHANIN2;
    input [10:0] TX_CHANIN3;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input TX_RESET;
    input TX_SERDES_REFCLK;
    input TX_SERDES_REFCLK_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module OBUFDS_GTE3 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTE3_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
    input [1:0] RXRECCLK_SEL;
endmodule

module OBUFDS_GTE4 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTE4_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
    input [1:0] RXRECCLK_SEL;
endmodule

module PCIE40E4 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AUTO_FLR_RESPONSE = "FALSE";
    parameter [1:0] AXISTEN_IF_CC_ALIGNMENT_MODE = 2'h0;
    parameter [23:0] AXISTEN_IF_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] AXISTEN_IF_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [1:0] AXISTEN_IF_CQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_CQ_EN_POISONED_MEM_WR = "FALSE";
    parameter AXISTEN_IF_ENABLE_256_TAGS = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE = "FALSE";
    parameter AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK = "TRUE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_EXT_512 = "FALSE";
    parameter AXISTEN_IF_EXT_512_CC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_CQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_LEGACY_MODE_ENABLE = "FALSE";
    parameter AXISTEN_IF_MSIX_FROM_RAM_PIPELINE = "FALSE";
    parameter AXISTEN_IF_MSIX_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_MSIX_TO_RAM_PIPELINE = "FALSE";
    parameter [1:0] AXISTEN_IF_RC_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter [1:0] AXISTEN_IF_RQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT = "FALSE";
    parameter AXISTEN_IF_TX_PARITY_EN = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CFG_BYPASS_MODE_ENABLE = "FALSE";
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter [15:0] DEBUG_AXI4ST_SPARE = 16'h0000;
    parameter [7:0] DEBUG_AXIST_DISABLE_FEATURE_BIT = 8'h00;
    parameter [3:0] DEBUG_CAR_SPARE = 4'h0;
    parameter [15:0] DEBUG_CFG_SPARE = 16'h0000;
    parameter [15:0] DEBUG_LL_SPARE = 16'h0000;
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW = "FALSE";
    parameter DEBUG_PL_DISABLE_SCRAMBLING = "FALSE";
    parameter DEBUG_PL_SIM_RESET_LFSR = "FALSE";
    parameter [15:0] DEBUG_PL_SPARE = 16'h0000;
    parameter DEBUG_TL_DISABLE_FC_TIMEOUT = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [15:0] DEBUG_TL_SPARE = 16'h0000;
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter DSN_CAP_ENABLE = "FALSE";
    parameter EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter HEADER_TYPE_OVERRIDE = "FALSE";
    parameter IS_SWITCH_PORT = "FALSE";
    parameter LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter LL_DISABLE_SCHED_TX_NAK = "FALSE";
    parameter LL_REPLAY_FROM_RAM_PIPELINE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter LL_REPLAY_TO_RAM_PIPELINE = "FALSE";
    parameter LL_RX_TLP_PARITY_GEN = "TRUE";
    parameter LL_TX_TLP_PARITY_CHK = "TRUE";
    parameter [15:0] LL_USER_SPARE = 16'h0000;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h250;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4 = 7;
    parameter [0:0] PF0_LINK_CONTROL_RCB = 1'h0;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [5:0] PF0_MSIX_VECTOR_COUNT = 6'h04;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter PL_CFG_STATE_ROBUSTNESS_ENABLE = "TRUE";
    parameter PL_DEEMPH_SOURCE_SELECT = "TRUE";
    parameter PL_DESKEW_ON_SKIP_IN_GEN12 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_LANE_REVERSAL = "FALSE";
    parameter [1:0] PL_DISABLE_LFSR_UPDATE_ON_SKP = 2'h0;
    parameter PL_DISABLE_RETRAIN_ON_EB_ERROR = "FALSE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter [15:0] PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR = 16'h0000;
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter [1:0] PL_EQ_ADAPT_DISABLE_COEFF_CHECK = 2'h0;
    parameter [1:0] PL_EQ_ADAPT_DISABLE_PRESET_CHECK = 2'h0;
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter [1:0] PL_EQ_BYPASS_PHASE23 = 2'h0;
    parameter [5:0] PL_EQ_DEFAULT_RX_PRESET_HINT = 6'h33;
    parameter [7:0] PL_EQ_DEFAULT_TX_PRESET = 8'h44;
    parameter PL_EQ_DISABLE_MISMATCH_CHECK = "TRUE";
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE0 = 2'h0;
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE1 = 2'h0;
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter PL_EQ_TX_8G_EQ_TS2_ENABLE = "FALSE";
    parameter PL_EXIT_LOOPBACK_ON_EI_ENTRY = "TRUE";
    parameter PL_INFER_EI_DISABLE_LPBK_ACTIVE = "TRUE";
    parameter PL_INFER_EI_DISABLE_REC_RC = "FALSE";
    parameter PL_INFER_EI_DISABLE_REC_SPD = "FALSE";
    parameter [31:0] PL_LANE0_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE10_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE11_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE12_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE13_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE14_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE15_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE1_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE2_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE3_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE4_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE5_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE6_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE7_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE8_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE9_EQ_CONTROL = 32'h00003F00;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_SPEED = 4'h4;
    parameter [4:0] PL_LINK_CAP_MAX_LINK_WIDTH = 5'h08;
    parameter integer PL_N_FTS = 255;
    parameter PL_QUIESCE_GUARANTEE_DISABLE = "FALSE";
    parameter PL_REDO_EQ_SOURCE_SELECT = "TRUE";
    parameter [7:0] PL_REPORT_ALL_PHY_ERRORS = 8'h00;
    parameter [1:0] PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN4 = 4'h0;
    parameter [1:0] PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN4 = 4'h0;
    parameter [1:0] PL_RX_L0S_EXIT_TO_RECOVERY = 2'h0;
    parameter [1:0] PL_SIM_FAST_LINK_TRAINING = 2'h0;
    parameter PL_SRIS_ENABLE = "FALSE";
    parameter [6:0] PL_SRIS_SKPOS_GEN_SPD_VEC = 7'h00;
    parameter [6:0] PL_SRIS_SKPOS_REC_SPD_VEC = 7'h00;
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PL_USER_SPARE = 16'h0000;
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h1500;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h003E8;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000100;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h00000;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0100;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter SPARE_BIT0 = "FALSE";
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter SPARE_BIT3 = "FALSE";
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter [3:0] SRIOV_CAP_ENABLE = 4'h0;
    parameter TL2CFG_IF_PARITY_CHK = "TRUE";
    parameter [1:0] TL_COMPLETION_RAM_NUM_TLPS = 2'h0;
    parameter [1:0] TL_COMPLETION_RAM_SIZE = 2'h1;
    parameter [11:0] TL_CREDITS_CD = 12'h000;
    parameter [7:0] TL_CREDITS_CH = 8'h00;
    parameter [11:0] TL_CREDITS_NPD = 12'h004;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h0E0;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TIME = 5'h02;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT = 5'h08;
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter [0:0] TL_POSTED_RAM_SIZE = 1'h0;
    parameter TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TL_TX_TLP_STRADDLE_ENABLE = "FALSE";
    parameter TL_TX_TLP_TERMINATE_PARITY = "FALSE";
    parameter [15:0] TL_USER_SPARE = 16'h0000;
    parameter TPH_FROM_RAM_PIPELINE = "FALSE";
    parameter TPH_TO_RAM_PIPELINE = "FALSE";
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h80;
    parameter [11:0] VFG0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    output [7:0] AXIUSEROUT;
    output [7:0] CFGBUSNUMBER;
    output [1:0] CFGCURRENTSPEED;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXVECPENDINGSTATUS;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output [4:0] CFGLOCALERROROUT;
    output CFGLOCALERRORVALID;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [1:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [12:0] CFGMSIXRAMADDRESS;
    output CFGMSIXRAMREADENABLE;
    output [3:0] CFGMSIXRAMWRITEBYTEENABLE;
    output [35:0] CFGMSIXRAMWRITEDATA;
    output [2:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [1:0] CFGRXPMSTATE;
    output [11:0] CFGTPHRAMADDRESS;
    output CFGTPHRAMREADENABLE;
    output [3:0] CFGTPHRAMWRITEBYTEENABLE;
    output [35:0] CFGTPHRAMWRITEDATA;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [1:0] CFGTXPMSTATE;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [31:0] DBGCTRL0OUT;
    output [31:0] DBGCTRL1OUT;
    output [255:0] DBGDATA0OUT;
    output [255:0] DBGDATA1OUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [87:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [8:0] MIREPLAYRAMADDRESS0;
    output [8:0] MIREPLAYRAMADDRESS1;
    output MIREPLAYRAMREADENABLE0;
    output MIREPLAYRAMREADENABLE1;
    output [127:0] MIREPLAYRAMWRITEDATA0;
    output [127:0] MIREPLAYRAMWRITEDATA1;
    output MIREPLAYRAMWRITEENABLE0;
    output MIREPLAYRAMWRITEENABLE1;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS1;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE0;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE1;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS1;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA0;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA1;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE0;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS1;
    output MIRXPOSTEDREQUESTRAMREADENABLE0;
    output MIRXPOSTEDREQUESTRAMREADENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS1;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA0;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA1;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE0;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE1;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [5:0] PCIERQSEQNUM0;
    output [5:0] PCIERQSEQNUM1;
    output PCIERQSEQNUMVLD0;
    output PCIERQSEQNUMVLD1;
    output [7:0] PCIERQTAG0;
    output [7:0] PCIERQTAG1;
    output [3:0] PCIERQTAGAV;
    output PCIERQTAGVLD0;
    output PCIERQTAGVLD1;
    output [3:0] PCIETFCNPDAV;
    output [3:0] PCIETFCNPHAV;
    output [1:0] PIPERX00EQCONTROL;
    output PIPERX00POLARITY;
    output [1:0] PIPERX01EQCONTROL;
    output PIPERX01POLARITY;
    output [1:0] PIPERX02EQCONTROL;
    output PIPERX02POLARITY;
    output [1:0] PIPERX03EQCONTROL;
    output PIPERX03POLARITY;
    output [1:0] PIPERX04EQCONTROL;
    output PIPERX04POLARITY;
    output [1:0] PIPERX05EQCONTROL;
    output PIPERX05POLARITY;
    output [1:0] PIPERX06EQCONTROL;
    output PIPERX06POLARITY;
    output [1:0] PIPERX07EQCONTROL;
    output PIPERX07POLARITY;
    output [1:0] PIPERX08EQCONTROL;
    output PIPERX08POLARITY;
    output [1:0] PIPERX09EQCONTROL;
    output PIPERX09POLARITY;
    output [1:0] PIPERX10EQCONTROL;
    output PIPERX10POLARITY;
    output [1:0] PIPERX11EQCONTROL;
    output PIPERX11POLARITY;
    output [1:0] PIPERX12EQCONTROL;
    output PIPERX12POLARITY;
    output [1:0] PIPERX13EQCONTROL;
    output PIPERX13POLARITY;
    output [1:0] PIPERX14EQCONTROL;
    output PIPERX14POLARITY;
    output [1:0] PIPERX15EQCONTROL;
    output PIPERX15POLARITY;
    output [5:0] PIPERXEQLPLFFS;
    output [3:0] PIPERXEQLPTXPRESET;
    output [1:0] PIPETX00CHARISK;
    output PIPETX00COMPLIANCE;
    output [31:0] PIPETX00DATA;
    output PIPETX00DATAVALID;
    output PIPETX00ELECIDLE;
    output [1:0] PIPETX00EQCONTROL;
    output [5:0] PIPETX00EQDEEMPH;
    output [1:0] PIPETX00POWERDOWN;
    output PIPETX00STARTBLOCK;
    output [1:0] PIPETX00SYNCHEADER;
    output [1:0] PIPETX01CHARISK;
    output PIPETX01COMPLIANCE;
    output [31:0] PIPETX01DATA;
    output PIPETX01DATAVALID;
    output PIPETX01ELECIDLE;
    output [1:0] PIPETX01EQCONTROL;
    output [5:0] PIPETX01EQDEEMPH;
    output [1:0] PIPETX01POWERDOWN;
    output PIPETX01STARTBLOCK;
    output [1:0] PIPETX01SYNCHEADER;
    output [1:0] PIPETX02CHARISK;
    output PIPETX02COMPLIANCE;
    output [31:0] PIPETX02DATA;
    output PIPETX02DATAVALID;
    output PIPETX02ELECIDLE;
    output [1:0] PIPETX02EQCONTROL;
    output [5:0] PIPETX02EQDEEMPH;
    output [1:0] PIPETX02POWERDOWN;
    output PIPETX02STARTBLOCK;
    output [1:0] PIPETX02SYNCHEADER;
    output [1:0] PIPETX03CHARISK;
    output PIPETX03COMPLIANCE;
    output [31:0] PIPETX03DATA;
    output PIPETX03DATAVALID;
    output PIPETX03ELECIDLE;
    output [1:0] PIPETX03EQCONTROL;
    output [5:0] PIPETX03EQDEEMPH;
    output [1:0] PIPETX03POWERDOWN;
    output PIPETX03STARTBLOCK;
    output [1:0] PIPETX03SYNCHEADER;
    output [1:0] PIPETX04CHARISK;
    output PIPETX04COMPLIANCE;
    output [31:0] PIPETX04DATA;
    output PIPETX04DATAVALID;
    output PIPETX04ELECIDLE;
    output [1:0] PIPETX04EQCONTROL;
    output [5:0] PIPETX04EQDEEMPH;
    output [1:0] PIPETX04POWERDOWN;
    output PIPETX04STARTBLOCK;
    output [1:0] PIPETX04SYNCHEADER;
    output [1:0] PIPETX05CHARISK;
    output PIPETX05COMPLIANCE;
    output [31:0] PIPETX05DATA;
    output PIPETX05DATAVALID;
    output PIPETX05ELECIDLE;
    output [1:0] PIPETX05EQCONTROL;
    output [5:0] PIPETX05EQDEEMPH;
    output [1:0] PIPETX05POWERDOWN;
    output PIPETX05STARTBLOCK;
    output [1:0] PIPETX05SYNCHEADER;
    output [1:0] PIPETX06CHARISK;
    output PIPETX06COMPLIANCE;
    output [31:0] PIPETX06DATA;
    output PIPETX06DATAVALID;
    output PIPETX06ELECIDLE;
    output [1:0] PIPETX06EQCONTROL;
    output [5:0] PIPETX06EQDEEMPH;
    output [1:0] PIPETX06POWERDOWN;
    output PIPETX06STARTBLOCK;
    output [1:0] PIPETX06SYNCHEADER;
    output [1:0] PIPETX07CHARISK;
    output PIPETX07COMPLIANCE;
    output [31:0] PIPETX07DATA;
    output PIPETX07DATAVALID;
    output PIPETX07ELECIDLE;
    output [1:0] PIPETX07EQCONTROL;
    output [5:0] PIPETX07EQDEEMPH;
    output [1:0] PIPETX07POWERDOWN;
    output PIPETX07STARTBLOCK;
    output [1:0] PIPETX07SYNCHEADER;
    output [1:0] PIPETX08CHARISK;
    output PIPETX08COMPLIANCE;
    output [31:0] PIPETX08DATA;
    output PIPETX08DATAVALID;
    output PIPETX08ELECIDLE;
    output [1:0] PIPETX08EQCONTROL;
    output [5:0] PIPETX08EQDEEMPH;
    output [1:0] PIPETX08POWERDOWN;
    output PIPETX08STARTBLOCK;
    output [1:0] PIPETX08SYNCHEADER;
    output [1:0] PIPETX09CHARISK;
    output PIPETX09COMPLIANCE;
    output [31:0] PIPETX09DATA;
    output PIPETX09DATAVALID;
    output PIPETX09ELECIDLE;
    output [1:0] PIPETX09EQCONTROL;
    output [5:0] PIPETX09EQDEEMPH;
    output [1:0] PIPETX09POWERDOWN;
    output PIPETX09STARTBLOCK;
    output [1:0] PIPETX09SYNCHEADER;
    output [1:0] PIPETX10CHARISK;
    output PIPETX10COMPLIANCE;
    output [31:0] PIPETX10DATA;
    output PIPETX10DATAVALID;
    output PIPETX10ELECIDLE;
    output [1:0] PIPETX10EQCONTROL;
    output [5:0] PIPETX10EQDEEMPH;
    output [1:0] PIPETX10POWERDOWN;
    output PIPETX10STARTBLOCK;
    output [1:0] PIPETX10SYNCHEADER;
    output [1:0] PIPETX11CHARISK;
    output PIPETX11COMPLIANCE;
    output [31:0] PIPETX11DATA;
    output PIPETX11DATAVALID;
    output PIPETX11ELECIDLE;
    output [1:0] PIPETX11EQCONTROL;
    output [5:0] PIPETX11EQDEEMPH;
    output [1:0] PIPETX11POWERDOWN;
    output PIPETX11STARTBLOCK;
    output [1:0] PIPETX11SYNCHEADER;
    output [1:0] PIPETX12CHARISK;
    output PIPETX12COMPLIANCE;
    output [31:0] PIPETX12DATA;
    output PIPETX12DATAVALID;
    output PIPETX12ELECIDLE;
    output [1:0] PIPETX12EQCONTROL;
    output [5:0] PIPETX12EQDEEMPH;
    output [1:0] PIPETX12POWERDOWN;
    output PIPETX12STARTBLOCK;
    output [1:0] PIPETX12SYNCHEADER;
    output [1:0] PIPETX13CHARISK;
    output PIPETX13COMPLIANCE;
    output [31:0] PIPETX13DATA;
    output PIPETX13DATAVALID;
    output PIPETX13ELECIDLE;
    output [1:0] PIPETX13EQCONTROL;
    output [5:0] PIPETX13EQDEEMPH;
    output [1:0] PIPETX13POWERDOWN;
    output PIPETX13STARTBLOCK;
    output [1:0] PIPETX13SYNCHEADER;
    output [1:0] PIPETX14CHARISK;
    output PIPETX14COMPLIANCE;
    output [31:0] PIPETX14DATA;
    output PIPETX14DATAVALID;
    output PIPETX14ELECIDLE;
    output [1:0] PIPETX14EQCONTROL;
    output [5:0] PIPETX14EQDEEMPH;
    output [1:0] PIPETX14POWERDOWN;
    output PIPETX14STARTBLOCK;
    output [1:0] PIPETX14SYNCHEADER;
    output [1:0] PIPETX15CHARISK;
    output PIPETX15COMPLIANCE;
    output [31:0] PIPETX15DATA;
    output PIPETX15DATAVALID;
    output PIPETX15ELECIDLE;
    output [1:0] PIPETX15EQCONTROL;
    output [5:0] PIPETX15EQDEEMPH;
    output [1:0] PIPETX15POWERDOWN;
    output PIPETX15STARTBLOCK;
    output [1:0] PIPETX15SYNCHEADER;
    output PIPETXDEEMPH;
    output [2:0] PIPETXMARGIN;
    output [1:0] PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PIPETXSWING;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output PLGEN34EQMISMATCH;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [31:0] USERSPAREOUT;
    input [7:0] AXIUSERIN;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVIDPF0;
    input [15:0] CFGDEVIDPF1;
    input [15:0] CFGDEVIDPF2;
    input [15:0] CFGDEVIDPF3;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [7:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [1:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [1:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [7:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [1:0] CFGINTERRUPTMSIXVECPENDING;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [9:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTDEBUGACCESS;
    input [7:0] CFGMGMTFUNCTIONNUMBER;
    input CFGMGMTREAD;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [35:0] CFGMSIXRAMREADDATA;
    input CFGPMASPML1ENTRYREJECT;
    input CFGPMASPMTXL0SENTRYDISABLE;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVIDPF0;
    input [7:0] CFGREVIDPF1;
    input [7:0] CFGREVIDPF2;
    input [7:0] CFGREVIDPF3;
    input [15:0] CFGSUBSYSIDPF0;
    input [15:0] CFGSUBSYSIDPF1;
    input [15:0] CFGSUBSYSIDPF2;
    input [15:0] CFGSUBSYSIDPF3;
    input [15:0] CFGSUBSYSVENDID;
    input [35:0] CFGTPHRAMREADDATA;
    input [15:0] CFGVENDID;
    input CFGVFFLRDONE;
    input [7:0] CFGVFFLRFUNCNUM;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKMIREPLAYRAM0;
    input CORECLKMIREPLAYRAM1;
    input CORECLKMIRXCOMPLETIONRAM0;
    input CORECLKMIRXCOMPLETIONRAM1;
    input CORECLKMIRXPOSTEDREQUESTRAM0;
    input CORECLKMIRXPOSTEDREQUESTRAM1;
    input [5:0] DBGSEL0;
    input [5:0] DBGSEL1;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [5:0] MIREPLAYRAMERRCOR;
    input [5:0] MIREPLAYRAMERRUNCOR;
    input [127:0] MIREPLAYRAMREADDATA0;
    input [127:0] MIREPLAYRAMREADDATA1;
    input [11:0] MIRXCOMPLETIONRAMERRCOR;
    input [11:0] MIRXCOMPLETIONRAMERRUNCOR;
    input [143:0] MIRXCOMPLETIONRAMREADDATA0;
    input [143:0] MIRXCOMPLETIONRAMREADDATA1;
    input [5:0] MIRXPOSTEDREQUESTRAMERRCOR;
    input [5:0] MIRXPOSTEDREQUESTRAMERRUNCOR;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA0;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA1;
    input [1:0] PCIECOMPLDELIVERED;
    input [7:0] PCIECOMPLDELIVEREDTAG0;
    input [7:0] PCIECOMPLDELIVEREDTAG1;
    input [1:0] PCIECQNPREQ;
    input PCIECQNPUSERCREDITRCVD;
    input PCIECQPIPELINEEMPTY;
    input PCIEPOSTEDREQDELIVERED;
    input PIPECLK;
    input PIPECLKEN;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX00CHARISK;
    input [31:0] PIPERX00DATA;
    input PIPERX00DATAVALID;
    input PIPERX00ELECIDLE;
    input PIPERX00EQDONE;
    input PIPERX00EQLPADAPTDONE;
    input PIPERX00EQLPLFFSSEL;
    input [17:0] PIPERX00EQLPNEWTXCOEFFORPRESET;
    input PIPERX00PHYSTATUS;
    input [1:0] PIPERX00STARTBLOCK;
    input [2:0] PIPERX00STATUS;
    input [1:0] PIPERX00SYNCHEADER;
    input PIPERX00VALID;
    input [1:0] PIPERX01CHARISK;
    input [31:0] PIPERX01DATA;
    input PIPERX01DATAVALID;
    input PIPERX01ELECIDLE;
    input PIPERX01EQDONE;
    input PIPERX01EQLPADAPTDONE;
    input PIPERX01EQLPLFFSSEL;
    input [17:0] PIPERX01EQLPNEWTXCOEFFORPRESET;
    input PIPERX01PHYSTATUS;
    input [1:0] PIPERX01STARTBLOCK;
    input [2:0] PIPERX01STATUS;
    input [1:0] PIPERX01SYNCHEADER;
    input PIPERX01VALID;
    input [1:0] PIPERX02CHARISK;
    input [31:0] PIPERX02DATA;
    input PIPERX02DATAVALID;
    input PIPERX02ELECIDLE;
    input PIPERX02EQDONE;
    input PIPERX02EQLPADAPTDONE;
    input PIPERX02EQLPLFFSSEL;
    input [17:0] PIPERX02EQLPNEWTXCOEFFORPRESET;
    input PIPERX02PHYSTATUS;
    input [1:0] PIPERX02STARTBLOCK;
    input [2:0] PIPERX02STATUS;
    input [1:0] PIPERX02SYNCHEADER;
    input PIPERX02VALID;
    input [1:0] PIPERX03CHARISK;
    input [31:0] PIPERX03DATA;
    input PIPERX03DATAVALID;
    input PIPERX03ELECIDLE;
    input PIPERX03EQDONE;
    input PIPERX03EQLPADAPTDONE;
    input PIPERX03EQLPLFFSSEL;
    input [17:0] PIPERX03EQLPNEWTXCOEFFORPRESET;
    input PIPERX03PHYSTATUS;
    input [1:0] PIPERX03STARTBLOCK;
    input [2:0] PIPERX03STATUS;
    input [1:0] PIPERX03SYNCHEADER;
    input PIPERX03VALID;
    input [1:0] PIPERX04CHARISK;
    input [31:0] PIPERX04DATA;
    input PIPERX04DATAVALID;
    input PIPERX04ELECIDLE;
    input PIPERX04EQDONE;
    input PIPERX04EQLPADAPTDONE;
    input PIPERX04EQLPLFFSSEL;
    input [17:0] PIPERX04EQLPNEWTXCOEFFORPRESET;
    input PIPERX04PHYSTATUS;
    input [1:0] PIPERX04STARTBLOCK;
    input [2:0] PIPERX04STATUS;
    input [1:0] PIPERX04SYNCHEADER;
    input PIPERX04VALID;
    input [1:0] PIPERX05CHARISK;
    input [31:0] PIPERX05DATA;
    input PIPERX05DATAVALID;
    input PIPERX05ELECIDLE;
    input PIPERX05EQDONE;
    input PIPERX05EQLPADAPTDONE;
    input PIPERX05EQLPLFFSSEL;
    input [17:0] PIPERX05EQLPNEWTXCOEFFORPRESET;
    input PIPERX05PHYSTATUS;
    input [1:0] PIPERX05STARTBLOCK;
    input [2:0] PIPERX05STATUS;
    input [1:0] PIPERX05SYNCHEADER;
    input PIPERX05VALID;
    input [1:0] PIPERX06CHARISK;
    input [31:0] PIPERX06DATA;
    input PIPERX06DATAVALID;
    input PIPERX06ELECIDLE;
    input PIPERX06EQDONE;
    input PIPERX06EQLPADAPTDONE;
    input PIPERX06EQLPLFFSSEL;
    input [17:0] PIPERX06EQLPNEWTXCOEFFORPRESET;
    input PIPERX06PHYSTATUS;
    input [1:0] PIPERX06STARTBLOCK;
    input [2:0] PIPERX06STATUS;
    input [1:0] PIPERX06SYNCHEADER;
    input PIPERX06VALID;
    input [1:0] PIPERX07CHARISK;
    input [31:0] PIPERX07DATA;
    input PIPERX07DATAVALID;
    input PIPERX07ELECIDLE;
    input PIPERX07EQDONE;
    input PIPERX07EQLPADAPTDONE;
    input PIPERX07EQLPLFFSSEL;
    input [17:0] PIPERX07EQLPNEWTXCOEFFORPRESET;
    input PIPERX07PHYSTATUS;
    input [1:0] PIPERX07STARTBLOCK;
    input [2:0] PIPERX07STATUS;
    input [1:0] PIPERX07SYNCHEADER;
    input PIPERX07VALID;
    input [1:0] PIPERX08CHARISK;
    input [31:0] PIPERX08DATA;
    input PIPERX08DATAVALID;
    input PIPERX08ELECIDLE;
    input PIPERX08EQDONE;
    input PIPERX08EQLPADAPTDONE;
    input PIPERX08EQLPLFFSSEL;
    input [17:0] PIPERX08EQLPNEWTXCOEFFORPRESET;
    input PIPERX08PHYSTATUS;
    input [1:0] PIPERX08STARTBLOCK;
    input [2:0] PIPERX08STATUS;
    input [1:0] PIPERX08SYNCHEADER;
    input PIPERX08VALID;
    input [1:0] PIPERX09CHARISK;
    input [31:0] PIPERX09DATA;
    input PIPERX09DATAVALID;
    input PIPERX09ELECIDLE;
    input PIPERX09EQDONE;
    input PIPERX09EQLPADAPTDONE;
    input PIPERX09EQLPLFFSSEL;
    input [17:0] PIPERX09EQLPNEWTXCOEFFORPRESET;
    input PIPERX09PHYSTATUS;
    input [1:0] PIPERX09STARTBLOCK;
    input [2:0] PIPERX09STATUS;
    input [1:0] PIPERX09SYNCHEADER;
    input PIPERX09VALID;
    input [1:0] PIPERX10CHARISK;
    input [31:0] PIPERX10DATA;
    input PIPERX10DATAVALID;
    input PIPERX10ELECIDLE;
    input PIPERX10EQDONE;
    input PIPERX10EQLPADAPTDONE;
    input PIPERX10EQLPLFFSSEL;
    input [17:0] PIPERX10EQLPNEWTXCOEFFORPRESET;
    input PIPERX10PHYSTATUS;
    input [1:0] PIPERX10STARTBLOCK;
    input [2:0] PIPERX10STATUS;
    input [1:0] PIPERX10SYNCHEADER;
    input PIPERX10VALID;
    input [1:0] PIPERX11CHARISK;
    input [31:0] PIPERX11DATA;
    input PIPERX11DATAVALID;
    input PIPERX11ELECIDLE;
    input PIPERX11EQDONE;
    input PIPERX11EQLPADAPTDONE;
    input PIPERX11EQLPLFFSSEL;
    input [17:0] PIPERX11EQLPNEWTXCOEFFORPRESET;
    input PIPERX11PHYSTATUS;
    input [1:0] PIPERX11STARTBLOCK;
    input [2:0] PIPERX11STATUS;
    input [1:0] PIPERX11SYNCHEADER;
    input PIPERX11VALID;
    input [1:0] PIPERX12CHARISK;
    input [31:0] PIPERX12DATA;
    input PIPERX12DATAVALID;
    input PIPERX12ELECIDLE;
    input PIPERX12EQDONE;
    input PIPERX12EQLPADAPTDONE;
    input PIPERX12EQLPLFFSSEL;
    input [17:0] PIPERX12EQLPNEWTXCOEFFORPRESET;
    input PIPERX12PHYSTATUS;
    input [1:0] PIPERX12STARTBLOCK;
    input [2:0] PIPERX12STATUS;
    input [1:0] PIPERX12SYNCHEADER;
    input PIPERX12VALID;
    input [1:0] PIPERX13CHARISK;
    input [31:0] PIPERX13DATA;
    input PIPERX13DATAVALID;
    input PIPERX13ELECIDLE;
    input PIPERX13EQDONE;
    input PIPERX13EQLPADAPTDONE;
    input PIPERX13EQLPLFFSSEL;
    input [17:0] PIPERX13EQLPNEWTXCOEFFORPRESET;
    input PIPERX13PHYSTATUS;
    input [1:0] PIPERX13STARTBLOCK;
    input [2:0] PIPERX13STATUS;
    input [1:0] PIPERX13SYNCHEADER;
    input PIPERX13VALID;
    input [1:0] PIPERX14CHARISK;
    input [31:0] PIPERX14DATA;
    input PIPERX14DATAVALID;
    input PIPERX14ELECIDLE;
    input PIPERX14EQDONE;
    input PIPERX14EQLPADAPTDONE;
    input PIPERX14EQLPLFFSSEL;
    input [17:0] PIPERX14EQLPNEWTXCOEFFORPRESET;
    input PIPERX14PHYSTATUS;
    input [1:0] PIPERX14STARTBLOCK;
    input [2:0] PIPERX14STATUS;
    input [1:0] PIPERX14SYNCHEADER;
    input PIPERX14VALID;
    input [1:0] PIPERX15CHARISK;
    input [31:0] PIPERX15DATA;
    input PIPERX15DATAVALID;
    input PIPERX15ELECIDLE;
    input PIPERX15EQDONE;
    input PIPERX15EQLPADAPTDONE;
    input PIPERX15EQLPLFFSSEL;
    input [17:0] PIPERX15EQLPNEWTXCOEFFORPRESET;
    input PIPERX15PHYSTATUS;
    input [1:0] PIPERX15STARTBLOCK;
    input [2:0] PIPERX15STATUS;
    input [1:0] PIPERX15SYNCHEADER;
    input PIPERX15VALID;
    input [17:0] PIPETX00EQCOEFF;
    input PIPETX00EQDONE;
    input [17:0] PIPETX01EQCOEFF;
    input PIPETX01EQDONE;
    input [17:0] PIPETX02EQCOEFF;
    input PIPETX02EQDONE;
    input [17:0] PIPETX03EQCOEFF;
    input PIPETX03EQDONE;
    input [17:0] PIPETX04EQCOEFF;
    input PIPETX04EQDONE;
    input [17:0] PIPETX05EQCOEFF;
    input PIPETX05EQDONE;
    input [17:0] PIPETX06EQCOEFF;
    input PIPETX06EQDONE;
    input [17:0] PIPETX07EQCOEFF;
    input PIPETX07EQDONE;
    input [17:0] PIPETX08EQCOEFF;
    input PIPETX08EQDONE;
    input [17:0] PIPETX09EQCOEFF;
    input PIPETX09EQDONE;
    input [17:0] PIPETX10EQCOEFF;
    input PIPETX10EQDONE;
    input [17:0] PIPETX11EQCOEFF;
    input PIPETX11EQDONE;
    input [17:0] PIPETX12EQCOEFF;
    input PIPETX12EQDONE;
    input [17:0] PIPETX13EQCOEFF;
    input PIPETX13EQDONE;
    input [17:0] PIPETX14EQCOEFF;
    input PIPETX14EQDONE;
    input [17:0] PIPETX15EQCOEFF;
    input PIPETX15EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input PLGEN34REDOEQSPEED;
    input PLGEN34REDOEQUALIZATION;
    input RESETN;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [61:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input USERCLK;
    input USERCLK2;
    input USERCLKEN;
    input [31:0] USERSPAREIN;
endmodule

module PCIE_3_1 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
    parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE = "FALSE";
    parameter DEBUG_PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF0_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_BIST_REGISTER = 8'h00;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter [15:0] PF0_DEVICE_ID = 16'h0000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF0_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
    parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF0_PB_CAP_VER = 4'h1;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter PF0_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF0_RBAR_NUM = 3'h1;
    parameter [7:0] PF0_REVISION_ID = 8'h00;
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF1_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_BIST_REGISTER = 8'h00;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [15:0] PF1_DEVICE_ID = 16'h0000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF1_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
    parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF1_PB_CAP_VER = 4'h1;
    parameter [7:0] PF1_PM_CAP_ID = 8'h01;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
    parameter PF1_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF1_RBAR_NUM = 3'h1;
    parameter [7:0] PF1_REVISION_ID = 8'h00;
    parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
    parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF1_TPHR_CAP_ENABLE = "FALSE";
    parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
    parameter PF2_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF2_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF2_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF2_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF2_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_BIST_REGISTER = 8'h00;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [15:0] PF2_DEVICE_ID = 16'h0000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF2_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF2_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF2_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF2_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF2_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF2_PB_CAP_NEXTPTR = 12'h000;
    parameter PF2_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF2_PB_CAP_VER = 4'h1;
    parameter [7:0] PF2_PM_CAP_ID = 8'h01;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF2_PM_CAP_VER_ID = 3'h3;
    parameter PF2_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF2_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF2_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF2_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF2_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF2_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF2_RBAR_NUM = 3'h1;
    parameter [7:0] PF2_REVISION_ID = 8'h00;
    parameter [4:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF2_SUBSYSTEM_ID = 16'h0000;
    parameter PF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF2_TPHR_CAP_ENABLE = "FALSE";
    parameter PF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF2_TPHR_CAP_VER = 4'h1;
    parameter PF3_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF3_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF3_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF3_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF3_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_BIST_REGISTER = 8'h00;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [15:0] PF3_DEVICE_ID = 16'h0000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF3_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF3_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF3_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF3_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF3_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF3_PB_CAP_NEXTPTR = 12'h000;
    parameter PF3_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF3_PB_CAP_VER = 4'h1;
    parameter [7:0] PF3_PM_CAP_ID = 8'h01;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF3_PM_CAP_VER_ID = 3'h3;
    parameter PF3_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF3_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF3_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF3_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF3_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF3_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF3_RBAR_NUM = 3'h1;
    parameter [7:0] PF3_REVISION_ID = 8'h00;
    parameter [4:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF3_SUBSYSTEM_ID = 16'h0000;
    parameter PF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF3_TPHR_CAP_ENABLE = "FALSE";
    parameter PF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF3_TPHR_CAP_VER = 4'h1;
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP = "TRUE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter PL_DISABLE_SCRAMBLING = "FALSE";
    parameter PL_DISABLE_SYNC_HEADER_FRAMING_ERROR = "FALSE";
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
    parameter [2:0] PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT = 3'h3;
    parameter [3:0] PL_EQ_DEFAULT_GEN3_TX_PRESET = 4'h4;
    parameter PL_EQ_PHASE01_RX_ADAPT = "FALSE";
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
    parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
    parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
    parameter integer PL_N_FTS_GEN1 = 255;
    parameter integer PL_N_FTS_GEN2 = 255;
    parameter integer PL_N_FTS_GEN3 = 255;
    parameter PL_REPORT_ALL_PHY_ERRORS = "TRUE";
    parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SRIOV_CAP_ENABLE = "FALSE";
    parameter TL_COMPLETION_RAM_SIZE_16K = "TRUE";
    parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [11:0] TL_CREDITS_CD = 12'h3E0;
    parameter [7:0] TL_CREDITS_CH = 8'h20;
    parameter [11:0] TL_CREDITS_NPD = 12'h028;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h198;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
    parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_MODE_ENABLE = "FALSE";
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TWO_LAYER_MODE_DLCMSM_ENABLE = "TRUE";
    parameter TWO_LAYER_MODE_ENABLE = "FALSE";
    parameter TWO_LAYER_MODE_WIDTH_256 = "TRUE";
    parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
    parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF0_PM_CAP_ID = 8'h01;
    parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
    parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF0_TPHR_CAP_ENABLE = "FALSE";
    parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF1_PM_CAP_ID = 8'h01;
    parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
    parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF1_TPHR_CAP_ENABLE = "FALSE";
    parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF2_PM_CAP_ID = 8'h01;
    parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
    parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF2_TPHR_CAP_ENABLE = "FALSE";
    parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF3_PM_CAP_ID = 8'h01;
    parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
    parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF3_TPHR_CAP_ENABLE = "FALSE";
    parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF4_PM_CAP_ID = 8'h01;
    parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
    parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF4_TPHR_CAP_ENABLE = "FALSE";
    parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF5_PM_CAP_ID = 8'h01;
    parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
    parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF5_TPHR_CAP_ENABLE = "FALSE";
    parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF6_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF6_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF6_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF6_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF6_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF6_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF6_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF6_PM_CAP_ID = 8'h01;
    parameter [7:0] VF6_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF6_PM_CAP_VER_ID = 3'h3;
    parameter VF6_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF6_TPHR_CAP_ENABLE = "FALSE";
    parameter VF6_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF6_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF6_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF6_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF6_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF6_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF7_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF7_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF7_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF7_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF7_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF7_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF7_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF7_PM_CAP_ID = 8'h01;
    parameter [7:0] VF7_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF7_PM_CAP_VER_ID = 3'h3;
    parameter VF7_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF7_TPHR_CAP_ENABLE = "FALSE";
    parameter VF7_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF7_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF7_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF7_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF7_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF7_TPHR_CAP_VER = 4'h1;
    output [2:0] CFGCURRENTSPEED;
    output [3:0] CFGDPASUBSTATECHANGE;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [7:0] CFGINTERRUPTMSIVFENABLE;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFAIL;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXSENT;
    output [7:0] CFGINTERRUPTMSIXVFENABLE;
    output [7:0] CFGINTERRUPTMSIXVFMASK;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output CFGLOCALERROR;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [2:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [3:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output [15:0] CFGPERFUNCSTATUSDATA;
    output CFGPERFUNCTIONUPDATEDONE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [3:0] CFGTPHFUNCTIONNUM;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [4:0] CFGTPHSTTADDRESS;
    output CFGTPHSTTREADENABLE;
    output [3:0] CFGTPHSTTWRITEBYTEVALID;
    output [31:0] CFGTPHSTTWRITEDATA;
    output CFGTPHSTTWRITEENABLE;
    output [7:0] CFGVFFLRINPROCESS;
    output [23:0] CFGVFPOWERSTATE;
    output [15:0] CFGVFSTATUS;
    output [7:0] CFGVFTPHREQUESTERENABLE;
    output [23:0] CFGVFTPHSTMODE;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [15:0] DBGDATAOUT;
    output DBGMCAPCSB;
    output [31:0] DBGMCAPDATA;
    output DBGMCAPEOS;
    output DBGMCAPERROR;
    output DBGMCAPMODE;
    output DBGMCAPRDATAVALID;
    output DBGMCAPRDWRB;
    output DBGMCAPRESET;
    output DBGPLDATABLOCKRECEIVEDAFTEREDS;
    output DBGPLGEN3FRAMINGERRORDETECTED;
    output DBGPLGEN3SYNCHEADERERRORDETECTED;
    output [7:0] DBGPLINFERREDRXELECTRICALIDLE;
    output [15:0] DRPDO;
    output DRPRDY;
    output LL2LMMASTERTLPSENT0;
    output LL2LMMASTERTLPSENT1;
    output [3:0] LL2LMMASTERTLPSENTTLPID0;
    output [3:0] LL2LMMASTERTLPSENTTLPID1;
    output [255:0] LL2LMMAXISRXTDATA;
    output [17:0] LL2LMMAXISRXTUSER;
    output [7:0] LL2LMMAXISRXTVALID;
    output [7:0] LL2LMSAXISTXTREADY;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [84:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [9:0] MICOMPLETIONRAMREADADDRESSAL;
    output [9:0] MICOMPLETIONRAMREADADDRESSAU;
    output [9:0] MICOMPLETIONRAMREADADDRESSBL;
    output [9:0] MICOMPLETIONRAMREADADDRESSBU;
    output [3:0] MICOMPLETIONRAMREADENABLEL;
    output [3:0] MICOMPLETIONRAMREADENABLEU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;
    output [71:0] MICOMPLETIONRAMWRITEDATAL;
    output [71:0] MICOMPLETIONRAMWRITEDATAU;
    output [3:0] MICOMPLETIONRAMWRITEENABLEL;
    output [3:0] MICOMPLETIONRAMWRITEENABLEU;
    output [8:0] MIREPLAYRAMADDRESS;
    output [1:0] MIREPLAYRAMREADENABLE;
    output [143:0] MIREPLAYRAMWRITEDATA;
    output [1:0] MIREPLAYRAMWRITEENABLE;
    output [8:0] MIREQUESTRAMREADADDRESSA;
    output [8:0] MIREQUESTRAMREADADDRESSB;
    output [3:0] MIREQUESTRAMREADENABLE;
    output [8:0] MIREQUESTRAMWRITEADDRESSA;
    output [8:0] MIREQUESTRAMWRITEADDRESSB;
    output [143:0] MIREQUESTRAMWRITEDATA;
    output [3:0] MIREQUESTRAMWRITEENABLE;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [3:0] PCIERQSEQNUM;
    output PCIERQSEQNUMVLD;
    output [5:0] PCIERQTAG;
    output [1:0] PCIERQTAGAV;
    output PCIERQTAGVLD;
    output [1:0] PCIETFCNPDAV;
    output [1:0] PCIETFCNPHAV;
    output [1:0] PIPERX0EQCONTROL;
    output [5:0] PIPERX0EQLPLFFS;
    output [3:0] PIPERX0EQLPTXPRESET;
    output [2:0] PIPERX0EQPRESET;
    output PIPERX0POLARITY;
    output [1:0] PIPERX1EQCONTROL;
    output [5:0] PIPERX1EQLPLFFS;
    output [3:0] PIPERX1EQLPTXPRESET;
    output [2:0] PIPERX1EQPRESET;
    output PIPERX1POLARITY;
    output [1:0] PIPERX2EQCONTROL;
    output [5:0] PIPERX2EQLPLFFS;
    output [3:0] PIPERX2EQLPTXPRESET;
    output [2:0] PIPERX2EQPRESET;
    output PIPERX2POLARITY;
    output [1:0] PIPERX3EQCONTROL;
    output [5:0] PIPERX3EQLPLFFS;
    output [3:0] PIPERX3EQLPTXPRESET;
    output [2:0] PIPERX3EQPRESET;
    output PIPERX3POLARITY;
    output [1:0] PIPERX4EQCONTROL;
    output [5:0] PIPERX4EQLPLFFS;
    output [3:0] PIPERX4EQLPTXPRESET;
    output [2:0] PIPERX4EQPRESET;
    output PIPERX4POLARITY;
    output [1:0] PIPERX5EQCONTROL;
    output [5:0] PIPERX5EQLPLFFS;
    output [3:0] PIPERX5EQLPTXPRESET;
    output [2:0] PIPERX5EQPRESET;
    output PIPERX5POLARITY;
    output [1:0] PIPERX6EQCONTROL;
    output [5:0] PIPERX6EQLPLFFS;
    output [3:0] PIPERX6EQLPTXPRESET;
    output [2:0] PIPERX6EQPRESET;
    output PIPERX6POLARITY;
    output [1:0] PIPERX7EQCONTROL;
    output [5:0] PIPERX7EQLPLFFS;
    output [3:0] PIPERX7EQLPTXPRESET;
    output [2:0] PIPERX7EQPRESET;
    output PIPERX7POLARITY;
    output [1:0] PIPETX0CHARISK;
    output PIPETX0COMPLIANCE;
    output [31:0] PIPETX0DATA;
    output PIPETX0DATAVALID;
    output PIPETX0DEEMPH;
    output PIPETX0ELECIDLE;
    output [1:0] PIPETX0EQCONTROL;
    output [5:0] PIPETX0EQDEEMPH;
    output [3:0] PIPETX0EQPRESET;
    output [2:0] PIPETX0MARGIN;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX0RATE;
    output PIPETX0RCVRDET;
    output PIPETX0RESET;
    output PIPETX0STARTBLOCK;
    output PIPETX0SWING;
    output [1:0] PIPETX0SYNCHEADER;
    output [1:0] PIPETX1CHARISK;
    output PIPETX1COMPLIANCE;
    output [31:0] PIPETX1DATA;
    output PIPETX1DATAVALID;
    output PIPETX1DEEMPH;
    output PIPETX1ELECIDLE;
    output [1:0] PIPETX1EQCONTROL;
    output [5:0] PIPETX1EQDEEMPH;
    output [3:0] PIPETX1EQPRESET;
    output [2:0] PIPETX1MARGIN;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX1RATE;
    output PIPETX1RCVRDET;
    output PIPETX1RESET;
    output PIPETX1STARTBLOCK;
    output PIPETX1SWING;
    output [1:0] PIPETX1SYNCHEADER;
    output [1:0] PIPETX2CHARISK;
    output PIPETX2COMPLIANCE;
    output [31:0] PIPETX2DATA;
    output PIPETX2DATAVALID;
    output PIPETX2DEEMPH;
    output PIPETX2ELECIDLE;
    output [1:0] PIPETX2EQCONTROL;
    output [5:0] PIPETX2EQDEEMPH;
    output [3:0] PIPETX2EQPRESET;
    output [2:0] PIPETX2MARGIN;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX2RATE;
    output PIPETX2RCVRDET;
    output PIPETX2RESET;
    output PIPETX2STARTBLOCK;
    output PIPETX2SWING;
    output [1:0] PIPETX2SYNCHEADER;
    output [1:0] PIPETX3CHARISK;
    output PIPETX3COMPLIANCE;
    output [31:0] PIPETX3DATA;
    output PIPETX3DATAVALID;
    output PIPETX3DEEMPH;
    output PIPETX3ELECIDLE;
    output [1:0] PIPETX3EQCONTROL;
    output [5:0] PIPETX3EQDEEMPH;
    output [3:0] PIPETX3EQPRESET;
    output [2:0] PIPETX3MARGIN;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX3RATE;
    output PIPETX3RCVRDET;
    output PIPETX3RESET;
    output PIPETX3STARTBLOCK;
    output PIPETX3SWING;
    output [1:0] PIPETX3SYNCHEADER;
    output [1:0] PIPETX4CHARISK;
    output PIPETX4COMPLIANCE;
    output [31:0] PIPETX4DATA;
    output PIPETX4DATAVALID;
    output PIPETX4DEEMPH;
    output PIPETX4ELECIDLE;
    output [1:0] PIPETX4EQCONTROL;
    output [5:0] PIPETX4EQDEEMPH;
    output [3:0] PIPETX4EQPRESET;
    output [2:0] PIPETX4MARGIN;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX4RATE;
    output PIPETX4RCVRDET;
    output PIPETX4RESET;
    output PIPETX4STARTBLOCK;
    output PIPETX4SWING;
    output [1:0] PIPETX4SYNCHEADER;
    output [1:0] PIPETX5CHARISK;
    output PIPETX5COMPLIANCE;
    output [31:0] PIPETX5DATA;
    output PIPETX5DATAVALID;
    output PIPETX5DEEMPH;
    output PIPETX5ELECIDLE;
    output [1:0] PIPETX5EQCONTROL;
    output [5:0] PIPETX5EQDEEMPH;
    output [3:0] PIPETX5EQPRESET;
    output [2:0] PIPETX5MARGIN;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX5RATE;
    output PIPETX5RCVRDET;
    output PIPETX5RESET;
    output PIPETX5STARTBLOCK;
    output PIPETX5SWING;
    output [1:0] PIPETX5SYNCHEADER;
    output [1:0] PIPETX6CHARISK;
    output PIPETX6COMPLIANCE;
    output [31:0] PIPETX6DATA;
    output PIPETX6DATAVALID;
    output PIPETX6DEEMPH;
    output PIPETX6ELECIDLE;
    output [1:0] PIPETX6EQCONTROL;
    output [5:0] PIPETX6EQDEEMPH;
    output [3:0] PIPETX6EQPRESET;
    output [2:0] PIPETX6MARGIN;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX6RATE;
    output PIPETX6RCVRDET;
    output PIPETX6RESET;
    output PIPETX6STARTBLOCK;
    output PIPETX6SWING;
    output [1:0] PIPETX6SYNCHEADER;
    output [1:0] PIPETX7CHARISK;
    output PIPETX7COMPLIANCE;
    output [31:0] PIPETX7DATA;
    output PIPETX7DATAVALID;
    output PIPETX7DEEMPH;
    output PIPETX7ELECIDLE;
    output [1:0] PIPETX7EQCONTROL;
    output [5:0] PIPETX7EQDEEMPH;
    output [3:0] PIPETX7EQPRESET;
    output [2:0] PIPETX7MARGIN;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PIPETX7RATE;
    output PIPETX7RCVRDET;
    output PIPETX7RESET;
    output PIPETX7STARTBLOCK;
    output PIPETX7SWING;
    output [1:0] PIPETX7SYNCHEADER;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [31:0] SPAREOUT;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVID;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [3:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [3:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [3:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [8:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [18:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTREAD;
    input CFGMGMTTYPE1CFGREGACCESS;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [2:0] CFGPERFUNCSTATUSCONTROL;
    input [3:0] CFGPERFUNCTIONNUMBER;
    input CFGPERFUNCTIONOUTPUTREQUEST;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [31:0] CFGTPHSTTREADDATA;
    input CFGTPHSTTREADDATAVALID;
    input [15:0] CFGVENDID;
    input [7:0] CFGVFFLRDONE;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKMICOMPLETIONRAML;
    input CORECLKMICOMPLETIONRAMU;
    input CORECLKMIREPLAYRAM;
    input CORECLKMIREQUESTRAM;
    input DBGCFGLOCALMGMTREGOVERRIDE;
    input [3:0] DBGDATASEL;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [13:0] LL2LMSAXISTXTUSER;
    input LL2LMSAXISTXTVALID;
    input [3:0] LL2LMTXTLPID0;
    input [3:0] LL2LMTXTLPID1;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [143:0] MICOMPLETIONRAMREADDATA;
    input [143:0] MIREPLAYRAMREADDATA;
    input [143:0] MIREQUESTRAMREADDATA;
    input PCIECQNPREQ;
    input PIPECLK;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX0CHARISK;
    input [31:0] PIPERX0DATA;
    input PIPERX0DATAVALID;
    input PIPERX0ELECIDLE;
    input PIPERX0EQDONE;
    input PIPERX0EQLPADAPTDONE;
    input PIPERX0EQLPLFFSSEL;
    input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
    input PIPERX0PHYSTATUS;
    input PIPERX0STARTBLOCK;
    input [2:0] PIPERX0STATUS;
    input [1:0] PIPERX0SYNCHEADER;
    input PIPERX0VALID;
    input [1:0] PIPERX1CHARISK;
    input [31:0] PIPERX1DATA;
    input PIPERX1DATAVALID;
    input PIPERX1ELECIDLE;
    input PIPERX1EQDONE;
    input PIPERX1EQLPADAPTDONE;
    input PIPERX1EQLPLFFSSEL;
    input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
    input PIPERX1PHYSTATUS;
    input PIPERX1STARTBLOCK;
    input [2:0] PIPERX1STATUS;
    input [1:0] PIPERX1SYNCHEADER;
    input PIPERX1VALID;
    input [1:0] PIPERX2CHARISK;
    input [31:0] PIPERX2DATA;
    input PIPERX2DATAVALID;
    input PIPERX2ELECIDLE;
    input PIPERX2EQDONE;
    input PIPERX2EQLPADAPTDONE;
    input PIPERX2EQLPLFFSSEL;
    input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
    input PIPERX2PHYSTATUS;
    input PIPERX2STARTBLOCK;
    input [2:0] PIPERX2STATUS;
    input [1:0] PIPERX2SYNCHEADER;
    input PIPERX2VALID;
    input [1:0] PIPERX3CHARISK;
    input [31:0] PIPERX3DATA;
    input PIPERX3DATAVALID;
    input PIPERX3ELECIDLE;
    input PIPERX3EQDONE;
    input PIPERX3EQLPADAPTDONE;
    input PIPERX3EQLPLFFSSEL;
    input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
    input PIPERX3PHYSTATUS;
    input PIPERX3STARTBLOCK;
    input [2:0] PIPERX3STATUS;
    input [1:0] PIPERX3SYNCHEADER;
    input PIPERX3VALID;
    input [1:0] PIPERX4CHARISK;
    input [31:0] PIPERX4DATA;
    input PIPERX4DATAVALID;
    input PIPERX4ELECIDLE;
    input PIPERX4EQDONE;
    input PIPERX4EQLPADAPTDONE;
    input PIPERX4EQLPLFFSSEL;
    input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
    input PIPERX4PHYSTATUS;
    input PIPERX4STARTBLOCK;
    input [2:0] PIPERX4STATUS;
    input [1:0] PIPERX4SYNCHEADER;
    input PIPERX4VALID;
    input [1:0] PIPERX5CHARISK;
    input [31:0] PIPERX5DATA;
    input PIPERX5DATAVALID;
    input PIPERX5ELECIDLE;
    input PIPERX5EQDONE;
    input PIPERX5EQLPADAPTDONE;
    input PIPERX5EQLPLFFSSEL;
    input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
    input PIPERX5PHYSTATUS;
    input PIPERX5STARTBLOCK;
    input [2:0] PIPERX5STATUS;
    input [1:0] PIPERX5SYNCHEADER;
    input PIPERX5VALID;
    input [1:0] PIPERX6CHARISK;
    input [31:0] PIPERX6DATA;
    input PIPERX6DATAVALID;
    input PIPERX6ELECIDLE;
    input PIPERX6EQDONE;
    input PIPERX6EQLPADAPTDONE;
    input PIPERX6EQLPLFFSSEL;
    input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
    input PIPERX6PHYSTATUS;
    input PIPERX6STARTBLOCK;
    input [2:0] PIPERX6STATUS;
    input [1:0] PIPERX6SYNCHEADER;
    input PIPERX6VALID;
    input [1:0] PIPERX7CHARISK;
    input [31:0] PIPERX7DATA;
    input PIPERX7DATAVALID;
    input PIPERX7ELECIDLE;
    input PIPERX7EQDONE;
    input PIPERX7EQLPADAPTDONE;
    input PIPERX7EQLPLFFSSEL;
    input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
    input PIPERX7PHYSTATUS;
    input PIPERX7STARTBLOCK;
    input [2:0] PIPERX7STATUS;
    input [1:0] PIPERX7SYNCHEADER;
    input PIPERX7VALID;
    input [17:0] PIPETX0EQCOEFF;
    input PIPETX0EQDONE;
    input [17:0] PIPETX1EQCOEFF;
    input PIPETX1EQDONE;
    input [17:0] PIPETX2EQCOEFF;
    input PIPETX2EQDONE;
    input [17:0] PIPETX3EQCOEFF;
    input PIPETX3EQDONE;
    input [17:0] PIPETX4EQCOEFF;
    input PIPETX4EQDONE;
    input [17:0] PIPETX5EQCOEFF;
    input PIPETX5EQDONE;
    input [17:0] PIPETX6EQCOEFF;
    input PIPETX6EQDONE;
    input [17:0] PIPETX7EQCOEFF;
    input PIPETX7EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input RESETN;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [59:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input [31:0] SPAREIN;
    input USERCLK;
endmodule

module SYSMONE1 (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter [15:0] INIT_58 = 16'h0;
    parameter [15:0] INIT_59 = 16'h0;
    parameter [15:0] INIT_5A = 16'h0;
    parameter [15:0] INIT_5B = 16'h0;
    parameter [15:0] INIT_5C = 16'h0;
    parameter [15:0] INIT_5D = 16'h0;
    parameter [15:0] INIT_5E = 16'h0;
    parameter [15:0] INIT_5F = 16'h0;
    parameter [15:0] INIT_60 = 16'h0;
    parameter [15:0] INIT_61 = 16'h0;
    parameter [15:0] INIT_62 = 16'h0;
    parameter [15:0] INIT_63 = 16'h0;
    parameter [15:0] INIT_64 = 16'h0;
    parameter [15:0] INIT_65 = 16'h0;
    parameter [15:0] INIT_66 = 16'h0;
    parameter [15:0] INIT_67 = 16'h0;
    parameter [15:0] INIT_68 = 16'h0;
    parameter [15:0] INIT_69 = 16'h0;
    parameter [15:0] INIT_6A = 16'h0;
    parameter [15:0] INIT_6B = 16'h0;
    parameter [15:0] INIT_6C = 16'h0;
    parameter [15:0] INIT_6D = 16'h0;
    parameter [15:0] INIT_6E = 16'h0;
    parameter [15:0] INIT_6F = 16'h0;
    parameter [15:0] INIT_70 = 16'h0;
    parameter [15:0] INIT_71 = 16'h0;
    parameter [15:0] INIT_72 = 16'h0;
    parameter [15:0] INIT_73 = 16'h0;
    parameter [15:0] INIT_74 = 16'h0;
    parameter [15:0] INIT_75 = 16'h0;
    parameter [15:0] INIT_76 = 16'h0;
    parameter [15:0] INIT_77 = 16'h0;
    parameter [15:0] INIT_78 = 16'h0;
    parameter [15:0] INIT_79 = 16'h0;
    parameter [15:0] INIT_7A = 16'h0;
    parameter [15:0] INIT_7B = 16'h0;
    parameter [15:0] INIT_7C = 16'h0;
    parameter [15:0] INIT_7D = 16'h0;
    parameter [15:0] INIT_7E = 16'h0;
    parameter [15:0] INIT_7F = 16'h0;
    parameter [0:0] IS_CONVSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DCLK_INVERTED = 1'b0;
    parameter SIM_MONITOR_FILE = "design.txt";
    parameter integer SYSMON_VUSER0_BANK = 0;
    parameter SYSMON_VUSER0_MONITOR = "NONE";
    parameter integer SYSMON_VUSER1_BANK = 0;
    parameter SYSMON_VUSER1_MONITOR = "NONE";
    parameter integer SYSMON_VUSER2_BANK = 0;
    parameter SYSMON_VUSER2_MONITOR = "NONE";
    parameter integer SYSMON_VUSER3_BANK = 0;
    parameter SYSMON_VUSER3_MONITOR = "NONE";
    output [15:0] ALM;
    output BUSY;
    output [5:0] CHANNEL;
    output [15:0] DO;
    output DRDY;
    output EOC;
    output EOS;
    output I2C_SCLK_TS;
    output I2C_SDA_TS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output [4:0] MUXADDR;
    output OT;
    input CONVST;
    input CONVSTCLK;
    input [7:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input I2C_SCLK;
    input I2C_SDA;
    input RESET;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input VN;
    input VP;
endmodule

module SYSMONE4 (...);
    parameter [15:0] COMMON_N_SOURCE = 16'hFFFF;
    parameter [15:0] INIT_40 = 16'h0000;
    parameter [15:0] INIT_41 = 16'h0000;
    parameter [15:0] INIT_42 = 16'h0000;
    parameter [15:0] INIT_43 = 16'h0000;
    parameter [15:0] INIT_44 = 16'h0000;
    parameter [15:0] INIT_45 = 16'h0000;
    parameter [15:0] INIT_46 = 16'h0000;
    parameter [15:0] INIT_47 = 16'h0000;
    parameter [15:0] INIT_48 = 16'h0000;
    parameter [15:0] INIT_49 = 16'h0000;
    parameter [15:0] INIT_4A = 16'h0000;
    parameter [15:0] INIT_4B = 16'h0000;
    parameter [15:0] INIT_4C = 16'h0000;
    parameter [15:0] INIT_4D = 16'h0000;
    parameter [15:0] INIT_4E = 16'h0000;
    parameter [15:0] INIT_4F = 16'h0000;
    parameter [15:0] INIT_50 = 16'h0000;
    parameter [15:0] INIT_51 = 16'h0000;
    parameter [15:0] INIT_52 = 16'h0000;
    parameter [15:0] INIT_53 = 16'h0000;
    parameter [15:0] INIT_54 = 16'h0000;
    parameter [15:0] INIT_55 = 16'h0000;
    parameter [15:0] INIT_56 = 16'h0000;
    parameter [15:0] INIT_57 = 16'h0000;
    parameter [15:0] INIT_58 = 16'h0000;
    parameter [15:0] INIT_59 = 16'h0000;
    parameter [15:0] INIT_5A = 16'h0000;
    parameter [15:0] INIT_5B = 16'h0000;
    parameter [15:0] INIT_5C = 16'h0000;
    parameter [15:0] INIT_5D = 16'h0000;
    parameter [15:0] INIT_5E = 16'h0000;
    parameter [15:0] INIT_5F = 16'h0000;
    parameter [15:0] INIT_60 = 16'h0000;
    parameter [15:0] INIT_61 = 16'h0000;
    parameter [15:0] INIT_62 = 16'h0000;
    parameter [15:0] INIT_63 = 16'h0000;
    parameter [15:0] INIT_64 = 16'h0000;
    parameter [15:0] INIT_65 = 16'h0000;
    parameter [15:0] INIT_66 = 16'h0000;
    parameter [15:0] INIT_67 = 16'h0000;
    parameter [15:0] INIT_68 = 16'h0000;
    parameter [15:0] INIT_69 = 16'h0000;
    parameter [15:0] INIT_6A = 16'h0000;
    parameter [15:0] INIT_6B = 16'h0000;
    parameter [15:0] INIT_6C = 16'h0000;
    parameter [15:0] INIT_6D = 16'h0000;
    parameter [15:0] INIT_6E = 16'h0000;
    parameter [15:0] INIT_6F = 16'h0000;
    parameter [15:0] INIT_70 = 16'h0000;
    parameter [15:0] INIT_71 = 16'h0000;
    parameter [15:0] INIT_72 = 16'h0000;
    parameter [15:0] INIT_73 = 16'h0000;
    parameter [15:0] INIT_74 = 16'h0000;
    parameter [15:0] INIT_75 = 16'h0000;
    parameter [15:0] INIT_76 = 16'h0000;
    parameter [15:0] INIT_77 = 16'h0000;
    parameter [15:0] INIT_78 = 16'h0000;
    parameter [15:0] INIT_79 = 16'h0000;
    parameter [15:0] INIT_7A = 16'h0000;
    parameter [15:0] INIT_7B = 16'h0000;
    parameter [15:0] INIT_7C = 16'h0000;
    parameter [15:0] INIT_7D = 16'h0000;
    parameter [15:0] INIT_7E = 16'h0000;
    parameter [15:0] INIT_7F = 16'h0000;
    parameter [0:0] IS_CONVSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DCLK_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MONITOR_FILE = "design.txt";
    parameter integer SYSMON_VUSER0_BANK = 0;
    parameter SYSMON_VUSER0_MONITOR = "NONE";
    parameter integer SYSMON_VUSER1_BANK = 0;
    parameter SYSMON_VUSER1_MONITOR = "NONE";
    parameter integer SYSMON_VUSER2_BANK = 0;
    parameter SYSMON_VUSER2_MONITOR = "NONE";
    parameter integer SYSMON_VUSER3_BANK = 0;
    parameter SYSMON_VUSER3_MONITOR = "NONE";
    output [15:0] ADC_DATA;
    output [15:0] ALM;
    output BUSY;
    output [5:0] CHANNEL;
    output [15:0] DO;
    output DRDY;
    output EOC;
    output EOS;
    output I2C_SCLK_TS;
    output I2C_SDA_TS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output [4:0] MUXADDR;
    output OT;
    output SMBALERT_TS;
    input CONVST;
    input CONVSTCLK;
    input [7:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input I2C_SCLK;
    input I2C_SDA;
    input RESET;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input VN;
    input VP;
endmodule

module DSP48E2 (...);
    parameter integer ACASCREG = 1;
    parameter integer ADREG = 1;
    parameter integer ALUMODEREG = 1;
    parameter AMULTSEL = "A";
    parameter integer AREG = 1;
    parameter AUTORESET_PATDET = "NO_RESET";
    parameter AUTORESET_PRIORITY = "RESET";
    parameter A_INPUT = "DIRECT";
    parameter integer BCASCREG = 1;
    parameter BMULTSEL = "B";
    parameter integer BREG = 1;
    parameter B_INPUT = "DIRECT";
    parameter integer CARRYINREG = 1;
    parameter integer CARRYINSELREG = 1;
    parameter integer CREG = 1;
    parameter integer DREG = 1;
    parameter integer INMODEREG = 1;
    parameter [3:0] IS_ALUMODE_INVERTED = 4'b0000;
    parameter [0:0] IS_CARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [4:0] IS_INMODE_INVERTED = 5'b00000;
    parameter [8:0] IS_OPMODE_INVERTED = 9'b000000000;
    parameter [0:0] IS_RSTALLCARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTALUMODE_INVERTED = 1'b0;
    parameter [0:0] IS_RSTA_INVERTED = 1'b0;
    parameter [0:0] IS_RSTB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTCTRL_INVERTED = 1'b0;
    parameter [0:0] IS_RSTC_INVERTED = 1'b0;
    parameter [0:0] IS_RSTD_INVERTED = 1'b0;
    parameter [0:0] IS_RSTINMODE_INVERTED = 1'b0;
    parameter [0:0] IS_RSTM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTP_INVERTED = 1'b0;
    parameter [47:0] MASK = 48'h3FFFFFFFFFFF;
    parameter integer MREG = 1;
    parameter integer OPMODEREG = 1;
    parameter [47:0] PATTERN = 48'h000000000000;
    parameter PREADDINSEL = "A";
    parameter integer PREG = 1;
    parameter [47:0] RND = 48'h000000000000;
    parameter SEL_MASK = "MASK";
    parameter SEL_PATTERN = "PATTERN";
    parameter USE_MULT = "MULTIPLY";
    parameter USE_PATTERN_DETECT = "NO_PATDET";
    parameter USE_SIMD = "ONE48";
    parameter USE_WIDEXOR = "FALSE";
    parameter XORSIMD = "XOR24_48_96";
    output [29:0] ACOUT;
    output [17:0] BCOUT;
    output CARRYCASCOUT;
    output [3:0] CARRYOUT;
    output MULTSIGNOUT;
    output OVERFLOW;
    output [47:0] P;
    output PATTERNBDETECT;
    output PATTERNDETECT;
    output [47:0] PCOUT;
    output UNDERFLOW;
    output [7:0] XOROUT;
    input [29:0] A;
    input [29:0] ACIN;
    input [3:0] ALUMODE;
    input [17:0] B;
    input [17:0] BCIN;
    input [47:0] C;
    input CARRYCASCIN;
    input CARRYIN;
    input [2:0] CARRYINSEL;
    input CEA1;
    input CEA2;
    input CEAD;
    input CEALUMODE;
    input CEB1;
    input CEB2;
    input CEC;
    input CECARRYIN;
    input CECTRL;
    input CED;
    input CEINMODE;
    input CEM;
    input CEP;
    (* clkbuf_sink *)
    input CLK;
    input [26:0] D;
    input [4:0] INMODE;
    input MULTSIGNIN;
    input [8:0] OPMODE;
    input [47:0] PCIN;
    input RSTA;
    input RSTALLCARRYIN;
    input RSTALUMODE;
    input RSTB;
    input RSTC;
    input RSTCTRL;
    input RSTD;
    input RSTINMODE;
    input RSTM;
    input RSTP;
endmodule

module FIFO18E2 (...);
    parameter CASCADE_ORDER = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter [35:0] INIT = 36'h000000000;
    parameter [0:0] IS_RDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RDEN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_WRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_WREN_INVERTED = 1'b0;
    parameter integer PROG_EMPTY_THRESH = 256;
    parameter integer PROG_FULL_THRESH = 256;
    parameter RDCOUNT_TYPE = "RAW_PNTR";
    parameter integer READ_WIDTH = 4;
    parameter REGISTER_MODE = "UNREGISTERED";
    parameter RSTREG_PRIORITY = "RSTREG";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [35:0] SRVAL = 36'h000000000;
    parameter WRCOUNT_TYPE = "RAW_PNTR";
    parameter integer WRITE_WIDTH = 4;
    output [31:0] CASDOUT;
    output [3:0] CASDOUTP;
    output CASNXTEMPTY;
    output CASPRVRDEN;
    output [31:0] DOUT;
    output [3:0] DOUTP;
    output EMPTY;
    output FULL;
    output PROGEMPTY;
    output PROGFULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output RDRSTBUSY;
    output [12:0] WRCOUNT;
    output WRERR;
    output WRRSTBUSY;
    input [31:0] CASDIN;
    input [3:0] CASDINP;
    input CASDOMUX;
    input CASDOMUXEN;
    input CASNXTRDEN;
    input CASOREGIMUX;
    input CASOREGIMUXEN;
    input CASPRVEMPTY;
    input [31:0] DIN;
    input [3:0] DINP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input REGCE;
    input RST;
    input RSTREG;
    input SLEEP;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module FIFO36E2 (...);
    parameter CASCADE_ORDER = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter EN_ECC_PIPE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter [71:0] INIT = 72'h000000000000000000;
    parameter [0:0] IS_RDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RDEN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_WRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_WREN_INVERTED = 1'b0;
    parameter integer PROG_EMPTY_THRESH = 256;
    parameter integer PROG_FULL_THRESH = 256;
    parameter RDCOUNT_TYPE = "RAW_PNTR";
    parameter integer READ_WIDTH = 4;
    parameter REGISTER_MODE = "UNREGISTERED";
    parameter RSTREG_PRIORITY = "RSTREG";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [71:0] SRVAL = 72'h000000000000000000;
    parameter WRCOUNT_TYPE = "RAW_PNTR";
    parameter integer WRITE_WIDTH = 4;
    output [63:0] CASDOUT;
    output [7:0] CASDOUTP;
    output CASNXTEMPTY;
    output CASPRVRDEN;
    output DBITERR;
    output [63:0] DOUT;
    output [7:0] DOUTP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output PROGEMPTY;
    output PROGFULL;
    output [13:0] RDCOUNT;
    output RDERR;
    output RDRSTBUSY;
    output SBITERR;
    output [13:0] WRCOUNT;
    output WRERR;
    output WRRSTBUSY;
    input [63:0] CASDIN;
    input [7:0] CASDINP;
    input CASDOMUX;
    input CASDOMUXEN;
    input CASNXTRDEN;
    input CASOREGIMUX;
    input CASOREGIMUXEN;
    input CASPRVEMPTY;
    input [63:0] DIN;
    input [7:0] DINP;
    input INJECTDBITERR;
    input INJECTSBITERR;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input REGCE;
    input RST;
    input RSTREG;
    input SLEEP;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module RAMB18E2 (...);
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter integer DOA_REG = 1;
    parameter integer DOB_REG = 1;
    parameter ENADDRENA = "FALSE";
    parameter ENADDRENB = "FALSE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [17:0] INIT_A = 18'h00000;
    parameter [17:0] INIT_B = 18'h00000;
    parameter INIT_FILE = "NONE";
    parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
    parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
    parameter RDADDRCHANGEA = "FALSE";
    parameter RDADDRCHANGEB = "FALSE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter RSTREG_PRIORITY_A = "RSTREG";
    parameter RSTREG_PRIORITY_B = "RSTREG";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [17:0] SRVAL_A = 18'h00000;
    parameter [17:0] SRVAL_B = 18'h00000;
    parameter WRITE_MODE_A = "NO_CHANGE";
    parameter WRITE_MODE_B = "NO_CHANGE";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [15:0] CASDOUTA;
    output [15:0] CASDOUTB;
    output [1:0] CASDOUTPA;
    output [1:0] CASDOUTPB;
    output [15:0] DOUTADOUT;
    output [15:0] DOUTBDOUT;
    output [1:0] DOUTPADOUTP;
    output [1:0] DOUTPBDOUTP;
    input [13:0] ADDRARDADDR;
    input [13:0] ADDRBWRADDR;
    input ADDRENA;
    input ADDRENB;
    input CASDIMUXA;
    input CASDIMUXB;
    input [15:0] CASDINA;
    input [15:0] CASDINB;
    input [1:0] CASDINPA;
    input [1:0] CASDINPB;
    input CASDOMUXA;
    input CASDOMUXB;
    input CASDOMUXEN_A;
    input CASDOMUXEN_B;
    input CASOREGIMUXA;
    input CASOREGIMUXB;
    input CASOREGIMUXEN_A;
    input CASOREGIMUXEN_B;
    (* clkbuf_sink *)
    input CLKARDCLK;
    (* clkbuf_sink *)
    input CLKBWRCLK;
    input [15:0] DINADIN;
    input [15:0] DINBDIN;
    input [1:0] DINPADINP;
    input [1:0] DINPBDINP;
    input ENARDEN;
    input ENBWREN;
    input REGCEAREGCE;
    input REGCEB;
    input RSTRAMARSTRAM;
    input RSTRAMB;
    input RSTREGARSTREG;
    input RSTREGB;
    input SLEEP;
    input [1:0] WEA;
    input [3:0] WEBWE;
endmodule

module RAMB36E2 (...);
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter integer DOA_REG = 1;
    parameter integer DOB_REG = 1;
    parameter ENADDRENA = "FALSE";
    parameter ENADDRENB = "FALSE";
    parameter EN_ECC_PIPE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [35:0] INIT_A = 36'h000000000;
    parameter [35:0] INIT_B = 36'h000000000;
    parameter INIT_FILE = "NONE";
    parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
    parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
    parameter RDADDRCHANGEA = "FALSE";
    parameter RDADDRCHANGEB = "FALSE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter RSTREG_PRIORITY_A = "RSTREG";
    parameter RSTREG_PRIORITY_B = "RSTREG";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [35:0] SRVAL_A = 36'h000000000;
    parameter [35:0] SRVAL_B = 36'h000000000;
    parameter WRITE_MODE_A = "NO_CHANGE";
    parameter WRITE_MODE_B = "NO_CHANGE";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [31:0] CASDOUTA;
    output [31:0] CASDOUTB;
    output [3:0] CASDOUTPA;
    output [3:0] CASDOUTPB;
    output CASOUTDBITERR;
    output CASOUTSBITERR;
    output DBITERR;
    output [31:0] DOUTADOUT;
    output [31:0] DOUTBDOUT;
    output [3:0] DOUTPADOUTP;
    output [3:0] DOUTPBDOUTP;
    output [7:0] ECCPARITY;
    output [8:0] RDADDRECC;
    output SBITERR;
    input [14:0] ADDRARDADDR;
    input [14:0] ADDRBWRADDR;
    input ADDRENA;
    input ADDRENB;
    input CASDIMUXA;
    input CASDIMUXB;
    input [31:0] CASDINA;
    input [31:0] CASDINB;
    input [3:0] CASDINPA;
    input [3:0] CASDINPB;
    input CASDOMUXA;
    input CASDOMUXB;
    input CASDOMUXEN_A;
    input CASDOMUXEN_B;
    input CASINDBITERR;
    input CASINSBITERR;
    input CASOREGIMUXA;
    input CASOREGIMUXB;
    input CASOREGIMUXEN_A;
    input CASOREGIMUXEN_B;
    (* clkbuf_sink *)
    input CLKARDCLK;
    (* clkbuf_sink *)
    input CLKBWRCLK;
    input [31:0] DINADIN;
    input [31:0] DINBDIN;
    input [3:0] DINPADINP;
    input [3:0] DINPBDINP;
    input ECCPIPECE;
    input ENARDEN;
    input ENBWREN;
    input INJECTDBITERR;
    input INJECTSBITERR;
    input REGCEAREGCE;
    input REGCEB;
    input RSTRAMARSTRAM;
    input RSTRAMB;
    input RSTREGARSTREG;
    input RSTREGB;
    input SLEEP;
    input [3:0] WEA;
    input [7:0] WEBWE;
endmodule

module URAM288 (...);
    parameter integer AUTO_SLEEP_LATENCY = 8;
    parameter integer AVG_CONS_INACTIVE_CYCLES = 10;
    parameter BWE_MODE_A = "PARITY_INTERLEAVED";
    parameter BWE_MODE_B = "PARITY_INTERLEAVED";
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter EN_AUTO_SLEEP_MODE = "FALSE";
    parameter EN_ECC_RD_A = "FALSE";
    parameter EN_ECC_RD_B = "FALSE";
    parameter EN_ECC_WR_A = "FALSE";
    parameter EN_ECC_WR_B = "FALSE";
    parameter IREG_PRE_A = "FALSE";
    parameter IREG_PRE_B = "FALSE";
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_EN_A_INVERTED = 1'b0;
    parameter [0:0] IS_EN_B_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_A_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_B_INVERTED = 1'b0;
    parameter [0:0] IS_RST_A_INVERTED = 1'b0;
    parameter [0:0] IS_RST_B_INVERTED = 1'b0;
    parameter MATRIX_ID = "NONE";
    parameter integer NUM_UNIQUE_SELF_ADDR_A = 1;
    parameter integer NUM_UNIQUE_SELF_ADDR_B = 1;
    parameter integer NUM_URAM_IN_MATRIX = 1;
    parameter OREG_A = "FALSE";
    parameter OREG_B = "FALSE";
    parameter OREG_ECC_A = "FALSE";
    parameter OREG_ECC_B = "FALSE";
    parameter REG_CAS_A = "FALSE";
    parameter REG_CAS_B = "FALSE";
    parameter RST_MODE_A = "SYNC";
    parameter RST_MODE_B = "SYNC";
    parameter [10:0] SELF_ADDR_A = 11'h000;
    parameter [10:0] SELF_ADDR_B = 11'h000;
    parameter [10:0] SELF_MASK_A = 11'h7FF;
    parameter [10:0] SELF_MASK_B = 11'h7FF;
    parameter USE_EXT_CE_A = "FALSE";
    parameter USE_EXT_CE_B = "FALSE";
    output [22:0] CAS_OUT_ADDR_A;
    output [22:0] CAS_OUT_ADDR_B;
    output [8:0] CAS_OUT_BWE_A;
    output [8:0] CAS_OUT_BWE_B;
    output CAS_OUT_DBITERR_A;
    output CAS_OUT_DBITERR_B;
    output [71:0] CAS_OUT_DIN_A;
    output [71:0] CAS_OUT_DIN_B;
    output [71:0] CAS_OUT_DOUT_A;
    output [71:0] CAS_OUT_DOUT_B;
    output CAS_OUT_EN_A;
    output CAS_OUT_EN_B;
    output CAS_OUT_RDACCESS_A;
    output CAS_OUT_RDACCESS_B;
    output CAS_OUT_RDB_WR_A;
    output CAS_OUT_RDB_WR_B;
    output CAS_OUT_SBITERR_A;
    output CAS_OUT_SBITERR_B;
    output DBITERR_A;
    output DBITERR_B;
    output [71:0] DOUT_A;
    output [71:0] DOUT_B;
    output RDACCESS_A;
    output RDACCESS_B;
    output SBITERR_A;
    output SBITERR_B;
    input [22:0] ADDR_A;
    input [22:0] ADDR_B;
    input [8:0] BWE_A;
    input [8:0] BWE_B;
    input [22:0] CAS_IN_ADDR_A;
    input [22:0] CAS_IN_ADDR_B;
    input [8:0] CAS_IN_BWE_A;
    input [8:0] CAS_IN_BWE_B;
    input CAS_IN_DBITERR_A;
    input CAS_IN_DBITERR_B;
    input [71:0] CAS_IN_DIN_A;
    input [71:0] CAS_IN_DIN_B;
    input [71:0] CAS_IN_DOUT_A;
    input [71:0] CAS_IN_DOUT_B;
    input CAS_IN_EN_A;
    input CAS_IN_EN_B;
    input CAS_IN_RDACCESS_A;
    input CAS_IN_RDACCESS_B;
    input CAS_IN_RDB_WR_A;
    input CAS_IN_RDB_WR_B;
    input CAS_IN_SBITERR_A;
    input CAS_IN_SBITERR_B;
    (* clkbuf_sink *)
    input CLK;
    input [71:0] DIN_A;
    input [71:0] DIN_B;
    input EN_A;
    input EN_B;
    input INJECT_DBITERR_A;
    input INJECT_DBITERR_B;
    input INJECT_SBITERR_A;
    input INJECT_SBITERR_B;
    input OREG_CE_A;
    input OREG_CE_B;
    input OREG_ECC_CE_A;
    input OREG_ECC_CE_B;
    input RDB_WR_A;
    input RDB_WR_B;
    input RST_A;
    input RST_B;
    input SLEEP;
endmodule

module URAM288_BASE (...);
    parameter integer AUTO_SLEEP_LATENCY = 8;
    parameter integer AVG_CONS_INACTIVE_CYCLES = 10;
    parameter BWE_MODE_A = "PARITY_INTERLEAVED";
    parameter BWE_MODE_B = "PARITY_INTERLEAVED";
    parameter EN_AUTO_SLEEP_MODE = "FALSE";
    parameter EN_ECC_RD_A = "FALSE";
    parameter EN_ECC_RD_B = "FALSE";
    parameter EN_ECC_WR_A = "FALSE";
    parameter EN_ECC_WR_B = "FALSE";
    parameter IREG_PRE_A = "FALSE";
    parameter IREG_PRE_B = "FALSE";
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_EN_A_INVERTED = 1'b0;
    parameter [0:0] IS_EN_B_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_A_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_B_INVERTED = 1'b0;
    parameter [0:0] IS_RST_A_INVERTED = 1'b0;
    parameter [0:0] IS_RST_B_INVERTED = 1'b0;
    parameter OREG_A = "FALSE";
    parameter OREG_B = "FALSE";
    parameter OREG_ECC_A = "FALSE";
    parameter OREG_ECC_B = "FALSE";
    parameter RST_MODE_A = "SYNC";
    parameter RST_MODE_B = "SYNC";
    parameter USE_EXT_CE_A = "FALSE";
    parameter USE_EXT_CE_B = "FALSE";
    output DBITERR_A;
    output DBITERR_B;
    output [71:0] DOUT_A;
    output [71:0] DOUT_B;
    output SBITERR_A;
    output SBITERR_B;
    input [22:0] ADDR_A;
    input [22:0] ADDR_B;
    input [8:0] BWE_A;
    input [8:0] BWE_B;
    (* clkbuf_sink *)
    input CLK;
    input [71:0] DIN_A;
    input [71:0] DIN_B;
    input EN_A;
    input EN_B;
    input INJECT_DBITERR_A;
    input INJECT_DBITERR_B;
    input INJECT_SBITERR_A;
    input INJECT_SBITERR_B;
    input OREG_CE_A;
    input OREG_CE_B;
    input OREG_ECC_CE_A;
    input OREG_ECC_CE_B;
    input RDB_WR_A;
    input RDB_WR_B;
    input RST_A;
    input RST_B;
    input SLEEP;
endmodule

module RAM128X1S (...);
    parameter [127:0] INIT = 128'h00000000000000000000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input A6;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM256X1D (...);
    parameter [255:0] INIT = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output DPO;
    output SPO;
    input [7:0] A;
    input D;
    input [7:0] DPRA;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM256X1S (...);
    parameter [255:0] INIT = 256'h0;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input [7:0] A;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32M (...);
    parameter [63:0] INIT_A = 64'h0000000000000000;
    parameter [63:0] INIT_B = 64'h0000000000000000;
    parameter [63:0] INIT_C = 64'h0000000000000000;
    parameter [63:0] INIT_D = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output [1:0] DOA;
    output [1:0] DOB;
    output [1:0] DOC;
    output [1:0] DOD;
    input [4:0] ADDRA;
    input [4:0] ADDRB;
    input [4:0] ADDRC;
    input [4:0] ADDRD;
    input [1:0] DIA;
    input [1:0] DIB;
    input [1:0] DIC;
    input [1:0] DID;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32M16 (...);
    parameter [63:0] INIT_A = 64'h0000000000000000;
    parameter [63:0] INIT_B = 64'h0000000000000000;
    parameter [63:0] INIT_C = 64'h0000000000000000;
    parameter [63:0] INIT_D = 64'h0000000000000000;
    parameter [63:0] INIT_E = 64'h0000000000000000;
    parameter [63:0] INIT_F = 64'h0000000000000000;
    parameter [63:0] INIT_G = 64'h0000000000000000;
    parameter [63:0] INIT_H = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output [1:0] DOA;
    output [1:0] DOB;
    output [1:0] DOC;
    output [1:0] DOD;
    output [1:0] DOE;
    output [1:0] DOF;
    output [1:0] DOG;
    output [1:0] DOH;
    input [4:0] ADDRA;
    input [4:0] ADDRB;
    input [4:0] ADDRC;
    input [4:0] ADDRD;
    input [4:0] ADDRE;
    input [4:0] ADDRF;
    input [4:0] ADDRG;
    input [4:0] ADDRH;
    input [1:0] DIA;
    input [1:0] DIB;
    input [1:0] DIC;
    input [1:0] DID;
    input [1:0] DIE;
    input [1:0] DIF;
    input [1:0] DIG;
    input [1:0] DIH;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32X1S (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM512X1S (...);
    parameter [511:0] INIT = 512'h0;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input [8:0] A;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64M (...);
    parameter [63:0] INIT_A = 64'h0000000000000000;
    parameter [63:0] INIT_B = 64'h0000000000000000;
    parameter [63:0] INIT_C = 64'h0000000000000000;
    parameter [63:0] INIT_D = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output DOA;
    output DOB;
    output DOC;
    output DOD;
    input [5:0] ADDRA;
    input [5:0] ADDRB;
    input [5:0] ADDRC;
    input [5:0] ADDRD;
    input DIA;
    input DIB;
    input DIC;
    input DID;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64M8 (...);
    parameter [63:0] INIT_A = 64'h0000000000000000;
    parameter [63:0] INIT_B = 64'h0000000000000000;
    parameter [63:0] INIT_C = 64'h0000000000000000;
    parameter [63:0] INIT_D = 64'h0000000000000000;
    parameter [63:0] INIT_E = 64'h0000000000000000;
    parameter [63:0] INIT_F = 64'h0000000000000000;
    parameter [63:0] INIT_G = 64'h0000000000000000;
    parameter [63:0] INIT_H = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output DOA;
    output DOB;
    output DOC;
    output DOD;
    output DOE;
    output DOF;
    output DOG;
    output DOH;
    input [5:0] ADDRA;
    input [5:0] ADDRB;
    input [5:0] ADDRC;
    input [5:0] ADDRD;
    input [5:0] ADDRE;
    input [5:0] ADDRF;
    input [5:0] ADDRG;
    input [5:0] ADDRH;
    input DIA;
    input DIB;
    input DIC;
    input DID;
    input DIE;
    input DIF;
    input DIG;
    input DIH;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64X1S (...);
    parameter [63:0] INIT = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module AND2B1L (...);
    parameter [0:0] IS_SRI_INVERTED = 1'b0;
    output O;
    input DI;
    input SRI;
endmodule

module CARRY8 (...);
    parameter CARRY_TYPE = "SINGLE_CY8";
    output [7:0] CO;
    output [7:0] O;
    input CI;
    input CI_TOP;
    input [7:0] DI;
    input [7:0] S;
endmodule

module CFGLUT5 (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    output CDO;
    output O5;
    output O6;
    input I4;
    input I3;
    input I2;
    input I1;
    input I0;
    input CDI;
    input CE;
    (* clkbuf_sink *)
    input CLK;
endmodule

module MUXF9 (...);
    output O;
    input I0;
    input I1;
    input S;
endmodule

module OR2L (...);
    parameter [0:0] IS_SRI_INVERTED = 1'b0;
    output O;
    input DI;
    input SRI;
endmodule

module BUFG_GT (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input CEMASK;
    input CLR;
    input CLRMASK;
    input [2:0] DIV;
    input I;
endmodule

module BUFG_GT_SYNC (...);
    output CESYNC;
    output CLRSYNC;
    input CE;
    input CLK;
    input CLR;
endmodule

module BUFG_PS (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFGCE (...);
    parameter CE_TYPE = "SYNC";
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    input CE;
    input I;
endmodule

module BUFGCE_1 (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input I;
endmodule

module BUFGCE_DIV (...);
    parameter integer BUFGCE_DIVIDE = 1;
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    input CE;
    input CLR;
    input I;
endmodule

module BUFGMUX (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_1 (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_CTRL (...);
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module MMCME3_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN2_INVERTED = 1'b0;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter STARTUP_WAIT = "FALSE";
    output CDDCDONE;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CDDCREQ;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input PWRDWN;
    input RST;
endmodule

module MMCME3_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module MMCME4_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN2_INVERTED = 1'b0;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 800.000;
    parameter STARTUP_WAIT = "FALSE";
    output CDDCDONE;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CDDCREQ;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input PWRDWN;
    input RST;
endmodule

module MMCME4_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module PLLE3_ADV (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 70.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter real CLKPFD_FREQ_MAX = 667.500;
    parameter real CLKPFD_FREQ_MIN = 70.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1335.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    input CLKFBIN;
    input CLKIN;
    input CLKOUTPHYEN;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PWRDWN;
    input RST;
endmodule

module PLLE3_BASE (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output LOCKED;
    input CLKFBIN;
    input CLKIN;
    input CLKOUTPHYEN;
    input PWRDWN;
    input RST;
endmodule

module PLLE4_ADV (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 70.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter real CLKPFD_FREQ_MAX = 667.500;
    parameter real CLKPFD_FREQ_MIN = 70.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1500.000;
    parameter real VCOCLK_FREQ_MIN = 750.000;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    input CLKFBIN;
    input CLKIN;
    input CLKOUTPHYEN;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PWRDWN;
    input RST;
endmodule

module PLLE4_BASE (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output LOCKED;
    input CLKFBIN;
    input CLKIN;
    input CLKOUTPHYEN;
    input PWRDWN;
    input RST;
endmodule

(* keep *)
module BSCANE2 (...);
    parameter DISABLE_JTAG = "FALSE";
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

module DNA_PORTE2 (...);
    parameter [95:0] SIM_DNA_VALUE = 96'h000000000000000000000000;
    output DOUT;
    input CLK;
    input DIN;
    input READ;
    input SHIFT;
endmodule

module EFUSE_USR (...);
    parameter [31:0] SIM_EFUSE_VALUE = 32'h00000000;
    output [31:0] EFUSEUSR;
endmodule

module FRAME_ECCE3 (...);
    output CRCERROR;
    output ECCERRORNOTSINGLE;
    output ECCERRORSINGLE;
    output ENDOFFRAME;
    output ENDOFSCAN;
    output [25:0] FAR;
    input [1:0] FARSEL;
    input ICAPBOTCLK;
    input ICAPTOPCLK;
endmodule

(* keep *)
module ICAPE3 (...);
    parameter [31:0] DEVICE_ID = 32'h03628093;
    parameter ICAP_AUTO_SWITCH = "DISABLE";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output AVAIL;
    output [31:0] O;
    output PRDONE;
    output PRERROR;
    input CLK;
    input CSIB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module MASTER_JTAG (...);
    output TDO;
    input TCK;
    input TDI;
    input TMS;
endmodule

(* keep *)
module STARTUPE3 (...);
    parameter PROG_USR = "FALSE";
    parameter real SIM_CCLK_FREQ = 0.0;
    output CFGCLK;
    output CFGMCLK;
    output [3:0] DI;
    output EOS;
    output PREQ;
    input [3:0] DO;
    input [3:0] DTS;
    input FCSBO;
    input FCSBTS;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

module USR_ACCESSE2 (...);
    output CFGCLK;
    output DATAVALID;
    output [31:0] DATA;
endmodule

(* keep *)
module BITSLICE_CONTROL (...);
    parameter CTRL_CLK = "EXTERNAL";
    parameter DIV_MODE = "DIV2";
    parameter EN_CLK_TO_EXT_NORTH = "DISABLE";
    parameter EN_CLK_TO_EXT_SOUTH = "DISABLE";
    parameter EN_DYN_ODLY_MODE = "FALSE";
    parameter EN_OTHER_NCLK = "FALSE";
    parameter EN_OTHER_PCLK = "FALSE";
    parameter IDLY_VT_TRACK = "TRUE";
    parameter INV_RXCLK = "FALSE";
    parameter ODLY_VT_TRACK = "TRUE";
    parameter QDLY_VT_TRACK = "TRUE";
    parameter [5:0] READ_IDLE_COUNT = 6'h00;
    parameter REFCLK_SRC = "PLLCLK";
    parameter integer ROUNDING_FACTOR = 16;
    parameter RXGATE_EXTEND = "FALSE";
    parameter RX_CLK_PHASE_N = "SHIFT_0";
    parameter RX_CLK_PHASE_P = "SHIFT_0";
    parameter RX_GATING = "DISABLE";
    parameter SELF_CALIBRATE = "ENABLE";
    parameter SERIAL_MODE = "FALSE";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter SIM_SPEEDUP = "FAST";
    parameter real SIM_VERSION = 2.0;
    parameter TX_GATING = "DISABLE";
    output CLK_TO_EXT_NORTH;
    output CLK_TO_EXT_SOUTH;
    output DLY_RDY;
    output [6:0] DYN_DCI;
    output NCLK_NIBBLE_OUT;
    output PCLK_NIBBLE_OUT;
    output [15:0] RIU_RD_DATA;
    output RIU_VALID;
    output [39:0] RX_BIT_CTRL_OUT0;
    output [39:0] RX_BIT_CTRL_OUT1;
    output [39:0] RX_BIT_CTRL_OUT2;
    output [39:0] RX_BIT_CTRL_OUT3;
    output [39:0] RX_BIT_CTRL_OUT4;
    output [39:0] RX_BIT_CTRL_OUT5;
    output [39:0] RX_BIT_CTRL_OUT6;
    output [39:0] TX_BIT_CTRL_OUT0;
    output [39:0] TX_BIT_CTRL_OUT1;
    output [39:0] TX_BIT_CTRL_OUT2;
    output [39:0] TX_BIT_CTRL_OUT3;
    output [39:0] TX_BIT_CTRL_OUT4;
    output [39:0] TX_BIT_CTRL_OUT5;
    output [39:0] TX_BIT_CTRL_OUT6;
    output [39:0] TX_BIT_CTRL_OUT_TRI;
    output VTC_RDY;
    input CLK_FROM_EXT;
    input EN_VTC;
    input NCLK_NIBBLE_IN;
    input PCLK_NIBBLE_IN;
    input [3:0] PHY_RDCS0;
    input [3:0] PHY_RDCS1;
    input [3:0] PHY_RDEN;
    input [3:0] PHY_WRCS0;
    input [3:0] PHY_WRCS1;
    input PLL_CLK;
    input REFCLK;
    input [5:0] RIU_ADDR;
    input RIU_CLK;
    input RIU_NIBBLE_SEL;
    input [15:0] RIU_WR_DATA;
    input RIU_WR_EN;
    input RST;
    input [39:0] RX_BIT_CTRL_IN0;
    input [39:0] RX_BIT_CTRL_IN1;
    input [39:0] RX_BIT_CTRL_IN2;
    input [39:0] RX_BIT_CTRL_IN3;
    input [39:0] RX_BIT_CTRL_IN4;
    input [39:0] RX_BIT_CTRL_IN5;
    input [39:0] RX_BIT_CTRL_IN6;
    input [3:0] TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN0;
    input [39:0] TX_BIT_CTRL_IN1;
    input [39:0] TX_BIT_CTRL_IN2;
    input [39:0] TX_BIT_CTRL_IN3;
    input [39:0] TX_BIT_CTRL_IN4;
    input [39:0] TX_BIT_CTRL_IN5;
    input [39:0] TX_BIT_CTRL_IN6;
    input [39:0] TX_BIT_CTRL_IN_TRI;
endmodule

(* keep *)
module DCIRESET (...);
    output LOCKED;
    input RST;
endmodule

module HPIO_VREF (...);
    parameter VREF_CNTR = "OFF";
    output VREF;
    input [6:0] FABRIC_VREF_TUNE;
endmodule

module IBUF_ANALOG (...);
    output O;
    (* iopad_external_pin *)
    input I;
endmodule

module IBUF_IBUFDISABLE (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
endmodule

module IBUF_INTERMDISABLE (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
endmodule

module IBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IFD_DELAY_VALUE = "AUTO";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_DIFF_OUT_IBUFDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
endmodule

module IBUFDS_DIFF_OUT_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input INTERMDISABLE;
endmodule

module IBUFDS_DPHY (...);
    parameter DIFF_TERM = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output HSRX_O;
    output LPRX_O_N;
    output LPRX_O_P;
    input HSRX_DISABLE;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input LPRX_DISABLE;
endmodule

module IBUFDS_IBUFDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
endmodule

module IBUFDS_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input INTERMDISABLE;
endmodule

module IBUFDSE3 (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input [3:0] OSC;
    input [1:0] OSC_EN;
endmodule

module IBUFE3 (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input OSC_EN;
    input VREF;
endmodule

(* keep *)
module IDELAYCTRL (...);
    parameter SIM_DEVICE = "7SERIES";
    output RDY;
    (* clkbuf_sink *)
    input REFCLK;
    input RST;
endmodule

module IDELAYE3 (...);
    parameter CASCADE = "NONE";
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_SRC = "IDATAIN";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter LOOPBACK = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output CASC_OUT;
    output [8:0] CNTVALUEOUT;
    output DATAOUT;
    input CASC_IN;
    input CASC_RETURN;
    input CE;
    (* clkbuf_sink *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input DATAIN;
    input EN_VTC;
    input IDATAIN;
    input INC;
    input LOAD;
    input RST;
endmodule

module IOBUF (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    output O;
    (* iopad_external_pin *)
    inout IO;
    input I;
    input T;
endmodule

module IOBUF_DCIEN (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input T;
endmodule

module IOBUF_INTERMDISABLE (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
    input T;
endmodule

module IOBUFDS (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    output O;
    (* iopad_external_pin *)
    inout IO;
    inout IOB;
    input I;
    input T;
endmodule

module IOBUFDS_DCIEN (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input T;
endmodule

module IOBUFDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input TM;
    input TS;
endmodule

module IOBUFDS_DIFF_OUT_DCIEN (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input TM;
    input TS;
endmodule

module IOBUFDS_DIFF_OUT_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
    input TM;
    input TS;
endmodule

module IOBUFDS_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
    input T;
endmodule

module IOBUFDSE3 (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    parameter USE_IBUFDISABLE = "FALSE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    inout IOB;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input [1:0] OSC_EN;
    input T;
endmodule

module IOBUFE3 (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    inout IO;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input OSC_EN;
    input T;
    input VREF;
endmodule

module ISERDESE3 (...);
    parameter integer DATA_WIDTH = 8;
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter FIFO_ENABLE = "FALSE";
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter IDDR_MODE = "FALSE";
    parameter [0:0] IS_CLK_B_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output FIFO_EMPTY;
    output INTERNAL_DIVCLK;
    output [7:0] Q;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    (* clkbuf_sink *)
    input CLK_B;
    input D;
    (* clkbuf_sink *)
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input RST;
endmodule

module KEEPER (...);
    inout O;
endmodule

module OBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
endmodule

module OBUFDS_DPHY (...);
    parameter IOSTANDARD = "DEFAULT";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input HSTX_I;
    input HSTX_T;
    input LPTX_I_N;
    input LPTX_I_P;
    input LPTX_T;
endmodule

module OBUFT (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter integer DRIVE = 12;
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    input I;
    input T;
endmodule

module OBUFTDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
    input T;
endmodule

module ODELAYE3 (...);
    parameter CASCADE = "NONE";
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output CASC_OUT;
    output [8:0] CNTVALUEOUT;
    output DATAOUT;
    input CASC_IN;
    input CASC_RETURN;
    input CE;
    (* clkbuf_sink *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input EN_VTC;
    input INC;
    input LOAD;
    input ODATAIN;
    input RST;
endmodule

module OSERDESE3 (...);
    parameter integer DATA_WIDTH = 8;
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter ODDR_MODE = "FALSE";
    parameter OSERDES_D_BYPASS = "FALSE";
    parameter OSERDES_T_BYPASS = "FALSE";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output OQ;
    output T_OUT;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    input [7:0] D;
    input RST;
    input T;
endmodule

module PULLDOWN (...);
    output O;
endmodule

module PULLUP (...);
    output O;
endmodule

module RIU_OR (...);
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output [15:0] RIU_RD_DATA;
    output RIU_RD_VALID;
    input [15:0] RIU_RD_DATA_LOW;
    input [15:0] RIU_RD_DATA_UPP;
    input RIU_RD_VALID_LOW;
    input RIU_RD_VALID_UPP;
endmodule

module RX_BITSLICE (...);
    parameter CASCADE = "TRUE";
    parameter DATA_TYPE = "NONE";
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter integer DELAY_VALUE_EXT = 0;
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter [0:0] IS_CLK_EXT_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_EXT_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    parameter UPDATE_MODE_EXT = "ASYNC";
    output [8:0] CNTVALUEOUT;
    output [8:0] CNTVALUEOUT_EXT;
    output FIFO_EMPTY;
    output FIFO_WRCLK_OUT;
    output [7:0] Q;
    output [39:0] RX_BIT_CTRL_OUT;
    output [39:0] TX_BIT_CTRL_OUT;
    input CE;
    input CE_EXT;
    input CLK;
    input CLK_EXT;
    input [8:0] CNTVALUEIN;
    input [8:0] CNTVALUEIN_EXT;
    input DATAIN;
    input EN_VTC;
    input EN_VTC_EXT;
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input INC;
    input INC_EXT;
    input LOAD;
    input LOAD_EXT;
    input RST;
    input RST_DLY;
    input RST_DLY_EXT;
    input [39:0] RX_BIT_CTRL_IN;
    input [39:0] TX_BIT_CTRL_IN;
endmodule

module RXTX_BITSLICE (...);
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_RX_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RX_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RX_RST_INVERTED = 1'b0;
    parameter [0:0] IS_TX_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_TX_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_TX_RST_INVERTED = 1'b0;
    parameter LOOPBACK = "FALSE";
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter ENABLE_PRE_EMPHASIS = "FALSE";
    parameter RX_DATA_TYPE = "NONE";
    parameter integer RX_DATA_WIDTH = 8;
    parameter RX_DELAY_FORMAT = "TIME";
    parameter RX_DELAY_TYPE = "FIXED";
    parameter integer RX_DELAY_VALUE = 0;
    parameter real RX_REFCLK_FREQUENCY = 300.0;
    parameter RX_UPDATE_MODE = "ASYNC";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter TBYTE_CTL = "TBYTE_IN";
    parameter integer TX_DATA_WIDTH = 8;
    parameter TX_DELAY_FORMAT = "TIME";
    parameter TX_DELAY_TYPE = "FIXED";
    parameter integer TX_DELAY_VALUE = 0;
    parameter TX_OUTPUT_PHASE_90 = "FALSE";
    parameter real TX_REFCLK_FREQUENCY = 300.0;
    parameter TX_UPDATE_MODE = "ASYNC";
    output FIFO_EMPTY;
    output FIFO_WRCLK_OUT;
    output O;
    output [7:0] Q;
    output [39:0] RX_BIT_CTRL_OUT;
    output [8:0] RX_CNTVALUEOUT;
    output [39:0] TX_BIT_CTRL_OUT;
    output [8:0] TX_CNTVALUEOUT;
    output T_OUT;
    input [7:0] D;
    input DATAIN;
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input [39:0] RX_BIT_CTRL_IN;
    input RX_CE;
    input RX_CLK;
    input [8:0] RX_CNTVALUEIN;
    input RX_EN_VTC;
    input RX_INC;
    input RX_LOAD;
    input RX_RST;
    input RX_RST_DLY;
    input T;
    input TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN;
    input TX_CE;
    input TX_CLK;
    input [8:0] TX_CNTVALUEIN;
    input TX_EN_VTC;
    input TX_INC;
    input TX_LOAD;
    input TX_RST;
    input TX_RST_DLY;
endmodule

module TX_BITSLICE (...);
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter ENABLE_PRE_EMPHASIS = "FALSE";
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter OUTPUT_PHASE_90 = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter TBYTE_CTL = "TBYTE_IN";
    parameter UPDATE_MODE = "ASYNC";
    output [8:0] CNTVALUEOUT;
    output O;
    output [39:0] RX_BIT_CTRL_OUT;
    output [39:0] TX_BIT_CTRL_OUT;
    output T_OUT;
    input CE;
    input CLK;
    input [8:0] CNTVALUEIN;
    input [7:0] D;
    input EN_VTC;
    input INC;
    input LOAD;
    input RST;
    input RST_DLY;
    input [39:0] RX_BIT_CTRL_IN;
    input T;
    input TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN;
endmodule

module TX_BITSLICE_TRI (...);
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter OUTPUT_PHASE_90 = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output [39:0] BIT_CTRL_OUT;
    output [8:0] CNTVALUEOUT;
    output TRI_OUT;
    input [39:0] BIT_CTRL_IN;
    input CE;
    input CLK;
    input [8:0] CNTVALUEIN;
    input EN_VTC;
    input INC;
    input LOAD;
    input RST;
    input RST_DLY;
endmodule

module HARD_SYNC (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter integer LATENCY = 2;
    output DOUT;
    (* clkbuf_sink *)
    input CLK;
    input DIN;
endmodule

module IDDRE1 (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter [0:0] IS_CB_INVERTED = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    input C;
    (* clkbuf_sink *)
    input CB;
    input D;
    input R;
endmodule

module LDCE (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_G_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    input CLR;
    input D;
    input G;
    input GE;
endmodule

module LDPE (...);
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_G_INVERTED = 1'b0;
    parameter [0:0] IS_PRE_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    input D;
    input G;
    input GE;
    input PRE;
endmodule

module ODDRE1 (...);
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter [0:0] SRVAL = 1'b0;
    output Q;
    (* clkbuf_sink *)
    input C;
    input D1;
    input D2;
    input SR;
endmodule

(* keep *)
module PS8 (...);
    output [7:0] ADMA2PLCACK;
    output [7:0] ADMA2PLTVLD;
    output DPAUDIOREFCLK;
    output DPAUXDATAOEN;
    output DPAUXDATAOUT;
    output DPLIVEVIDEODEOUT;
    output [31:0] DPMAXISMIXEDAUDIOTDATA;
    output DPMAXISMIXEDAUDIOTID;
    output DPMAXISMIXEDAUDIOTVALID;
    output DPSAXISAUDIOTREADY;
    output DPVIDEOOUTHSYNC;
    output [35:0] DPVIDEOOUTPIXEL1;
    output DPVIDEOOUTVSYNC;
    output DPVIDEOREFCLK;
    output EMIOCAN0PHYTX;
    output EMIOCAN1PHYTX;
    output [1:0] EMIOENET0DMABUSWIDTH;
    output EMIOENET0DMATXENDTOG;
    output [93:0] EMIOENET0GEMTSUTIMERCNT;
    output [7:0] EMIOENET0GMIITXD;
    output EMIOENET0GMIITXEN;
    output EMIOENET0GMIITXER;
    output EMIOENET0MDIOMDC;
    output EMIOENET0MDIOO;
    output EMIOENET0MDIOTN;
    output [7:0] EMIOENET0RXWDATA;
    output EMIOENET0RXWEOP;
    output EMIOENET0RXWERR;
    output EMIOENET0RXWFLUSH;
    output EMIOENET0RXWSOP;
    output [44:0] EMIOENET0RXWSTATUS;
    output EMIOENET0RXWWR;
    output [2:0] EMIOENET0SPEEDMODE;
    output EMIOENET0TXRRD;
    output [3:0] EMIOENET0TXRSTATUS;
    output [1:0] EMIOENET1DMABUSWIDTH;
    output EMIOENET1DMATXENDTOG;
    output [7:0] EMIOENET1GMIITXD;
    output EMIOENET1GMIITXEN;
    output EMIOENET1GMIITXER;
    output EMIOENET1MDIOMDC;
    output EMIOENET1MDIOO;
    output EMIOENET1MDIOTN;
    output [7:0] EMIOENET1RXWDATA;
    output EMIOENET1RXWEOP;
    output EMIOENET1RXWERR;
    output EMIOENET1RXWFLUSH;
    output EMIOENET1RXWSOP;
    output [44:0] EMIOENET1RXWSTATUS;
    output EMIOENET1RXWWR;
    output [2:0] EMIOENET1SPEEDMODE;
    output EMIOENET1TXRRD;
    output [3:0] EMIOENET1TXRSTATUS;
    output [1:0] EMIOENET2DMABUSWIDTH;
    output EMIOENET2DMATXENDTOG;
    output [7:0] EMIOENET2GMIITXD;
    output EMIOENET2GMIITXEN;
    output EMIOENET2GMIITXER;
    output EMIOENET2MDIOMDC;
    output EMIOENET2MDIOO;
    output EMIOENET2MDIOTN;
    output [7:0] EMIOENET2RXWDATA;
    output EMIOENET2RXWEOP;
    output EMIOENET2RXWERR;
    output EMIOENET2RXWFLUSH;
    output EMIOENET2RXWSOP;
    output [44:0] EMIOENET2RXWSTATUS;
    output EMIOENET2RXWWR;
    output [2:0] EMIOENET2SPEEDMODE;
    output EMIOENET2TXRRD;
    output [3:0] EMIOENET2TXRSTATUS;
    output [1:0] EMIOENET3DMABUSWIDTH;
    output EMIOENET3DMATXENDTOG;
    output [7:0] EMIOENET3GMIITXD;
    output EMIOENET3GMIITXEN;
    output EMIOENET3GMIITXER;
    output EMIOENET3MDIOMDC;
    output EMIOENET3MDIOO;
    output EMIOENET3MDIOTN;
    output [7:0] EMIOENET3RXWDATA;
    output EMIOENET3RXWEOP;
    output EMIOENET3RXWERR;
    output EMIOENET3RXWFLUSH;
    output EMIOENET3RXWSOP;
    output [44:0] EMIOENET3RXWSTATUS;
    output EMIOENET3RXWWR;
    output [2:0] EMIOENET3SPEEDMODE;
    output EMIOENET3TXRRD;
    output [3:0] EMIOENET3TXRSTATUS;
    output EMIOGEM0DELAYREQRX;
    output EMIOGEM0DELAYREQTX;
    output EMIOGEM0PDELAYREQRX;
    output EMIOGEM0PDELAYREQTX;
    output EMIOGEM0PDELAYRESPRX;
    output EMIOGEM0PDELAYRESPTX;
    output EMIOGEM0RXSOF;
    output EMIOGEM0SYNCFRAMERX;
    output EMIOGEM0SYNCFRAMETX;
    output EMIOGEM0TSUTIMERCMPVAL;
    output EMIOGEM0TXRFIXEDLAT;
    output EMIOGEM0TXSOF;
    output EMIOGEM1DELAYREQRX;
    output EMIOGEM1DELAYREQTX;
    output EMIOGEM1PDELAYREQRX;
    output EMIOGEM1PDELAYREQTX;
    output EMIOGEM1PDELAYRESPRX;
    output EMIOGEM1PDELAYRESPTX;
    output EMIOGEM1RXSOF;
    output EMIOGEM1SYNCFRAMERX;
    output EMIOGEM1SYNCFRAMETX;
    output EMIOGEM1TSUTIMERCMPVAL;
    output EMIOGEM1TXRFIXEDLAT;
    output EMIOGEM1TXSOF;
    output EMIOGEM2DELAYREQRX;
    output EMIOGEM2DELAYREQTX;
    output EMIOGEM2PDELAYREQRX;
    output EMIOGEM2PDELAYREQTX;
    output EMIOGEM2PDELAYRESPRX;
    output EMIOGEM2PDELAYRESPTX;
    output EMIOGEM2RXSOF;
    output EMIOGEM2SYNCFRAMERX;
    output EMIOGEM2SYNCFRAMETX;
    output EMIOGEM2TSUTIMERCMPVAL;
    output EMIOGEM2TXRFIXEDLAT;
    output EMIOGEM2TXSOF;
    output EMIOGEM3DELAYREQRX;
    output EMIOGEM3DELAYREQTX;
    output EMIOGEM3PDELAYREQRX;
    output EMIOGEM3PDELAYREQTX;
    output EMIOGEM3PDELAYRESPRX;
    output EMIOGEM3PDELAYRESPTX;
    output EMIOGEM3RXSOF;
    output EMIOGEM3SYNCFRAMERX;
    output EMIOGEM3SYNCFRAMETX;
    output EMIOGEM3TSUTIMERCMPVAL;
    output EMIOGEM3TXRFIXEDLAT;
    output EMIOGEM3TXSOF;
    output [95:0] EMIOGPIOO;
    output [95:0] EMIOGPIOTN;
    output EMIOI2C0SCLO;
    output EMIOI2C0SCLTN;
    output EMIOI2C0SDAO;
    output EMIOI2C0SDATN;
    output EMIOI2C1SCLO;
    output EMIOI2C1SCLTN;
    output EMIOI2C1SDAO;
    output EMIOI2C1SDATN;
    output EMIOSDIO0BUSPOWER;
    output [2:0] EMIOSDIO0BUSVOLT;
    output EMIOSDIO0CLKOUT;
    output EMIOSDIO0CMDENA;
    output EMIOSDIO0CMDOUT;
    output [7:0] EMIOSDIO0DATAENA;
    output [7:0] EMIOSDIO0DATAOUT;
    output EMIOSDIO0LEDCONTROL;
    output EMIOSDIO1BUSPOWER;
    output [2:0] EMIOSDIO1BUSVOLT;
    output EMIOSDIO1CLKOUT;
    output EMIOSDIO1CMDENA;
    output EMIOSDIO1CMDOUT;
    output [7:0] EMIOSDIO1DATAENA;
    output [7:0] EMIOSDIO1DATAOUT;
    output EMIOSDIO1LEDCONTROL;
    output EMIOSPI0MO;
    output EMIOSPI0MOTN;
    output EMIOSPI0SCLKO;
    output EMIOSPI0SCLKTN;
    output EMIOSPI0SO;
    output EMIOSPI0SSNTN;
    output [2:0] EMIOSPI0SSON;
    output EMIOSPI0STN;
    output EMIOSPI1MO;
    output EMIOSPI1MOTN;
    output EMIOSPI1SCLKO;
    output EMIOSPI1SCLKTN;
    output EMIOSPI1SO;
    output EMIOSPI1SSNTN;
    output [2:0] EMIOSPI1SSON;
    output EMIOSPI1STN;
    output [2:0] EMIOTTC0WAVEO;
    output [2:0] EMIOTTC1WAVEO;
    output [2:0] EMIOTTC2WAVEO;
    output [2:0] EMIOTTC3WAVEO;
    output EMIOU2DSPORTVBUSCTRLUSB30;
    output EMIOU2DSPORTVBUSCTRLUSB31;
    output EMIOU3DSPORTVBUSCTRLUSB30;
    output EMIOU3DSPORTVBUSCTRLUSB31;
    output EMIOUART0DTRN;
    output EMIOUART0RTSN;
    output EMIOUART0TX;
    output EMIOUART1DTRN;
    output EMIOUART1RTSN;
    output EMIOUART1TX;
    output EMIOWDT0RSTO;
    output EMIOWDT1RSTO;
    output FMIOGEM0FIFORXCLKTOPLBUFG;
    output FMIOGEM0FIFOTXCLKTOPLBUFG;
    output FMIOGEM1FIFORXCLKTOPLBUFG;
    output FMIOGEM1FIFOTXCLKTOPLBUFG;
    output FMIOGEM2FIFORXCLKTOPLBUFG;
    output FMIOGEM2FIFOTXCLKTOPLBUFG;
    output FMIOGEM3FIFORXCLKTOPLBUFG;
    output FMIOGEM3FIFOTXCLKTOPLBUFG;
    output FMIOGEMTSUCLKTOPLBUFG;
    output [31:0] FTMGPO;
    output [7:0] GDMA2PLCACK;
    output [7:0] GDMA2PLTVLD;
    output [39:0] MAXIGP0ARADDR;
    output [1:0] MAXIGP0ARBURST;
    output [3:0] MAXIGP0ARCACHE;
    output [15:0] MAXIGP0ARID;
    output [7:0] MAXIGP0ARLEN;
    output MAXIGP0ARLOCK;
    output [2:0] MAXIGP0ARPROT;
    output [3:0] MAXIGP0ARQOS;
    output [2:0] MAXIGP0ARSIZE;
    output [15:0] MAXIGP0ARUSER;
    output MAXIGP0ARVALID;
    output [39:0] MAXIGP0AWADDR;
    output [1:0] MAXIGP0AWBURST;
    output [3:0] MAXIGP0AWCACHE;
    output [15:0] MAXIGP0AWID;
    output [7:0] MAXIGP0AWLEN;
    output MAXIGP0AWLOCK;
    output [2:0] MAXIGP0AWPROT;
    output [3:0] MAXIGP0AWQOS;
    output [2:0] MAXIGP0AWSIZE;
    output [15:0] MAXIGP0AWUSER;
    output MAXIGP0AWVALID;
    output MAXIGP0BREADY;
    output MAXIGP0RREADY;
    output [127:0] MAXIGP0WDATA;
    output MAXIGP0WLAST;
    output [15:0] MAXIGP0WSTRB;
    output MAXIGP0WVALID;
    output [39:0] MAXIGP1ARADDR;
    output [1:0] MAXIGP1ARBURST;
    output [3:0] MAXIGP1ARCACHE;
    output [15:0] MAXIGP1ARID;
    output [7:0] MAXIGP1ARLEN;
    output MAXIGP1ARLOCK;
    output [2:0] MAXIGP1ARPROT;
    output [3:0] MAXIGP1ARQOS;
    output [2:0] MAXIGP1ARSIZE;
    output [15:0] MAXIGP1ARUSER;
    output MAXIGP1ARVALID;
    output [39:0] MAXIGP1AWADDR;
    output [1:0] MAXIGP1AWBURST;
    output [3:0] MAXIGP1AWCACHE;
    output [15:0] MAXIGP1AWID;
    output [7:0] MAXIGP1AWLEN;
    output MAXIGP1AWLOCK;
    output [2:0] MAXIGP1AWPROT;
    output [3:0] MAXIGP1AWQOS;
    output [2:0] MAXIGP1AWSIZE;
    output [15:0] MAXIGP1AWUSER;
    output MAXIGP1AWVALID;
    output MAXIGP1BREADY;
    output MAXIGP1RREADY;
    output [127:0] MAXIGP1WDATA;
    output MAXIGP1WLAST;
    output [15:0] MAXIGP1WSTRB;
    output MAXIGP1WVALID;
    output [39:0] MAXIGP2ARADDR;
    output [1:0] MAXIGP2ARBURST;
    output [3:0] MAXIGP2ARCACHE;
    output [15:0] MAXIGP2ARID;
    output [7:0] MAXIGP2ARLEN;
    output MAXIGP2ARLOCK;
    output [2:0] MAXIGP2ARPROT;
    output [3:0] MAXIGP2ARQOS;
    output [2:0] MAXIGP2ARSIZE;
    output [15:0] MAXIGP2ARUSER;
    output MAXIGP2ARVALID;
    output [39:0] MAXIGP2AWADDR;
    output [1:0] MAXIGP2AWBURST;
    output [3:0] MAXIGP2AWCACHE;
    output [15:0] MAXIGP2AWID;
    output [7:0] MAXIGP2AWLEN;
    output MAXIGP2AWLOCK;
    output [2:0] MAXIGP2AWPROT;
    output [3:0] MAXIGP2AWQOS;
    output [2:0] MAXIGP2AWSIZE;
    output [15:0] MAXIGP2AWUSER;
    output MAXIGP2AWVALID;
    output MAXIGP2BREADY;
    output MAXIGP2RREADY;
    output [127:0] MAXIGP2WDATA;
    output MAXIGP2WLAST;
    output [15:0] MAXIGP2WSTRB;
    output MAXIGP2WVALID;
    output OSCRTCCLK;
    output [3:0] PLCLK;
    output PMUAIBAFIFMFPDREQ;
    output PMUAIBAFIFMLPDREQ;
    output [46:0] PMUERRORTOPL;
    output [31:0] PMUPLGPO;
    output PSPLEVENTO;
    output [63:0] PSPLIRQFPD;
    output [99:0] PSPLIRQLPD;
    output [3:0] PSPLSTANDBYWFE;
    output [3:0] PSPLSTANDBYWFI;
    output PSPLTRACECTL;
    output [31:0] PSPLTRACEDATA;
    output [3:0] PSPLTRIGACK;
    output [3:0] PSPLTRIGGER;
    output PSS_ALTO_CORE_PAD_MGTTXN0OUT;
    output PSS_ALTO_CORE_PAD_MGTTXN1OUT;
    output PSS_ALTO_CORE_PAD_MGTTXN2OUT;
    output PSS_ALTO_CORE_PAD_MGTTXN3OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP0OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP1OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP2OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP3OUT;
    output PSS_ALTO_CORE_PAD_PADO;
    output RPUEVENTO0;
    output RPUEVENTO1;
    output [43:0] SACEFPDACADDR;
    output [2:0] SACEFPDACPROT;
    output [3:0] SACEFPDACSNOOP;
    output SACEFPDACVALID;
    output SACEFPDARREADY;
    output SACEFPDAWREADY;
    output [5:0] SACEFPDBID;
    output [1:0] SACEFPDBRESP;
    output SACEFPDBUSER;
    output SACEFPDBVALID;
    output SACEFPDCDREADY;
    output SACEFPDCRREADY;
    output [127:0] SACEFPDRDATA;
    output [5:0] SACEFPDRID;
    output SACEFPDRLAST;
    output [3:0] SACEFPDRRESP;
    output SACEFPDRUSER;
    output SACEFPDRVALID;
    output SACEFPDWREADY;
    output SAXIACPARREADY;
    output SAXIACPAWREADY;
    output [4:0] SAXIACPBID;
    output [1:0] SAXIACPBRESP;
    output SAXIACPBVALID;
    output [127:0] SAXIACPRDATA;
    output [4:0] SAXIACPRID;
    output SAXIACPRLAST;
    output [1:0] SAXIACPRRESP;
    output SAXIACPRVALID;
    output SAXIACPWREADY;
    output SAXIGP0ARREADY;
    output SAXIGP0AWREADY;
    output [5:0] SAXIGP0BID;
    output [1:0] SAXIGP0BRESP;
    output SAXIGP0BVALID;
    output [3:0] SAXIGP0RACOUNT;
    output [7:0] SAXIGP0RCOUNT;
    output [127:0] SAXIGP0RDATA;
    output [5:0] SAXIGP0RID;
    output SAXIGP0RLAST;
    output [1:0] SAXIGP0RRESP;
    output SAXIGP0RVALID;
    output [3:0] SAXIGP0WACOUNT;
    output [7:0] SAXIGP0WCOUNT;
    output SAXIGP0WREADY;
    output SAXIGP1ARREADY;
    output SAXIGP1AWREADY;
    output [5:0] SAXIGP1BID;
    output [1:0] SAXIGP1BRESP;
    output SAXIGP1BVALID;
    output [3:0] SAXIGP1RACOUNT;
    output [7:0] SAXIGP1RCOUNT;
    output [127:0] SAXIGP1RDATA;
    output [5:0] SAXIGP1RID;
    output SAXIGP1RLAST;
    output [1:0] SAXIGP1RRESP;
    output SAXIGP1RVALID;
    output [3:0] SAXIGP1WACOUNT;
    output [7:0] SAXIGP1WCOUNT;
    output SAXIGP1WREADY;
    output SAXIGP2ARREADY;
    output SAXIGP2AWREADY;
    output [5:0] SAXIGP2BID;
    output [1:0] SAXIGP2BRESP;
    output SAXIGP2BVALID;
    output [3:0] SAXIGP2RACOUNT;
    output [7:0] SAXIGP2RCOUNT;
    output [127:0] SAXIGP2RDATA;
    output [5:0] SAXIGP2RID;
    output SAXIGP2RLAST;
    output [1:0] SAXIGP2RRESP;
    output SAXIGP2RVALID;
    output [3:0] SAXIGP2WACOUNT;
    output [7:0] SAXIGP2WCOUNT;
    output SAXIGP2WREADY;
    output SAXIGP3ARREADY;
    output SAXIGP3AWREADY;
    output [5:0] SAXIGP3BID;
    output [1:0] SAXIGP3BRESP;
    output SAXIGP3BVALID;
    output [3:0] SAXIGP3RACOUNT;
    output [7:0] SAXIGP3RCOUNT;
    output [127:0] SAXIGP3RDATA;
    output [5:0] SAXIGP3RID;
    output SAXIGP3RLAST;
    output [1:0] SAXIGP3RRESP;
    output SAXIGP3RVALID;
    output [3:0] SAXIGP3WACOUNT;
    output [7:0] SAXIGP3WCOUNT;
    output SAXIGP3WREADY;
    output SAXIGP4ARREADY;
    output SAXIGP4AWREADY;
    output [5:0] SAXIGP4BID;
    output [1:0] SAXIGP4BRESP;
    output SAXIGP4BVALID;
    output [3:0] SAXIGP4RACOUNT;
    output [7:0] SAXIGP4RCOUNT;
    output [127:0] SAXIGP4RDATA;
    output [5:0] SAXIGP4RID;
    output SAXIGP4RLAST;
    output [1:0] SAXIGP4RRESP;
    output SAXIGP4RVALID;
    output [3:0] SAXIGP4WACOUNT;
    output [7:0] SAXIGP4WCOUNT;
    output SAXIGP4WREADY;
    output SAXIGP5ARREADY;
    output SAXIGP5AWREADY;
    output [5:0] SAXIGP5BID;
    output [1:0] SAXIGP5BRESP;
    output SAXIGP5BVALID;
    output [3:0] SAXIGP5RACOUNT;
    output [7:0] SAXIGP5RCOUNT;
    output [127:0] SAXIGP5RDATA;
    output [5:0] SAXIGP5RID;
    output SAXIGP5RLAST;
    output [1:0] SAXIGP5RRESP;
    output SAXIGP5RVALID;
    output [3:0] SAXIGP5WACOUNT;
    output [7:0] SAXIGP5WCOUNT;
    output SAXIGP5WREADY;
    output SAXIGP6ARREADY;
    output SAXIGP6AWREADY;
    output [5:0] SAXIGP6BID;
    output [1:0] SAXIGP6BRESP;
    output SAXIGP6BVALID;
    output [3:0] SAXIGP6RACOUNT;
    output [7:0] SAXIGP6RCOUNT;
    output [127:0] SAXIGP6RDATA;
    output [5:0] SAXIGP6RID;
    output SAXIGP6RLAST;
    output [1:0] SAXIGP6RRESP;
    output SAXIGP6RVALID;
    output [3:0] SAXIGP6WACOUNT;
    output [7:0] SAXIGP6WCOUNT;
    output SAXIGP6WREADY;
    inout [3:0] PSS_ALTO_CORE_PAD_BOOTMODE;
    inout PSS_ALTO_CORE_PAD_CLK;
    inout PSS_ALTO_CORE_PAD_DONEB;
    inout [17:0] PSS_ALTO_CORE_PAD_DRAMA;
    inout PSS_ALTO_CORE_PAD_DRAMACTN;
    inout PSS_ALTO_CORE_PAD_DRAMALERTN;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMBA;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMBG;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCK;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCKE;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCKN;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCSN;
    inout [8:0] PSS_ALTO_CORE_PAD_DRAMDM;
    inout [71:0] PSS_ALTO_CORE_PAD_DRAMDQ;
    inout [8:0] PSS_ALTO_CORE_PAD_DRAMDQS;
    inout [8:0] PSS_ALTO_CORE_PAD_DRAMDQSN;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMODT;
    inout PSS_ALTO_CORE_PAD_DRAMPARITY;
    inout PSS_ALTO_CORE_PAD_DRAMRAMRSTN;
    inout PSS_ALTO_CORE_PAD_ERROROUT;
    inout PSS_ALTO_CORE_PAD_ERRORSTATUS;
    inout PSS_ALTO_CORE_PAD_INITB;
    inout PSS_ALTO_CORE_PAD_JTAGTCK;
    inout PSS_ALTO_CORE_PAD_JTAGTDI;
    inout PSS_ALTO_CORE_PAD_JTAGTDO;
    inout PSS_ALTO_CORE_PAD_JTAGTMS;
    inout [77:0] PSS_ALTO_CORE_PAD_MIO;
    inout PSS_ALTO_CORE_PAD_PORB;
    inout PSS_ALTO_CORE_PAD_PROGB;
    inout PSS_ALTO_CORE_PAD_RCALIBINOUT;
    inout PSS_ALTO_CORE_PAD_SRSTB;
    inout PSS_ALTO_CORE_PAD_ZQ;
    input [7:0] ADMAFCICLK;
    input AIBPMUAFIFMFPDACK;
    input AIBPMUAFIFMLPDACK;
    input DDRCEXTREFRESHRANK0REQ;
    input DDRCEXTREFRESHRANK1REQ;
    input DDRCREFRESHPLCLK;
    input DPAUXDATAIN;
    input DPEXTERNALCUSTOMEVENT1;
    input DPEXTERNALCUSTOMEVENT2;
    input DPEXTERNALVSYNCEVENT;
    input DPHOTPLUGDETECT;
    input [7:0] DPLIVEGFXALPHAIN;
    input [35:0] DPLIVEGFXPIXEL1IN;
    input DPLIVEVIDEOINDE;
    input DPLIVEVIDEOINHSYNC;
    input [35:0] DPLIVEVIDEOINPIXEL1;
    input DPLIVEVIDEOINVSYNC;
    input DPMAXISMIXEDAUDIOTREADY;
    input DPSAXISAUDIOCLK;
    input [31:0] DPSAXISAUDIOTDATA;
    input DPSAXISAUDIOTID;
    input DPSAXISAUDIOTVALID;
    input DPVIDEOINCLK;
    input EMIOCAN0PHYRX;
    input EMIOCAN1PHYRX;
    input EMIOENET0DMATXSTATUSTOG;
    input EMIOENET0EXTINTIN;
    input EMIOENET0GMIICOL;
    input EMIOENET0GMIICRS;
    input EMIOENET0GMIIRXCLK;
    input [7:0] EMIOENET0GMIIRXD;
    input EMIOENET0GMIIRXDV;
    input EMIOENET0GMIIRXER;
    input EMIOENET0GMIITXCLK;
    input EMIOENET0MDIOI;
    input EMIOENET0RXWOVERFLOW;
    input EMIOENET0TXRCONTROL;
    input [7:0] EMIOENET0TXRDATA;
    input EMIOENET0TXRDATARDY;
    input EMIOENET0TXREOP;
    input EMIOENET0TXRERR;
    input EMIOENET0TXRFLUSHED;
    input EMIOENET0TXRSOP;
    input EMIOENET0TXRUNDERFLOW;
    input EMIOENET0TXRVALID;
    input EMIOENET1DMATXSTATUSTOG;
    input EMIOENET1EXTINTIN;
    input EMIOENET1GMIICOL;
    input EMIOENET1GMIICRS;
    input EMIOENET1GMIIRXCLK;
    input [7:0] EMIOENET1GMIIRXD;
    input EMIOENET1GMIIRXDV;
    input EMIOENET1GMIIRXER;
    input EMIOENET1GMIITXCLK;
    input EMIOENET1MDIOI;
    input EMIOENET1RXWOVERFLOW;
    input EMIOENET1TXRCONTROL;
    input [7:0] EMIOENET1TXRDATA;
    input EMIOENET1TXRDATARDY;
    input EMIOENET1TXREOP;
    input EMIOENET1TXRERR;
    input EMIOENET1TXRFLUSHED;
    input EMIOENET1TXRSOP;
    input EMIOENET1TXRUNDERFLOW;
    input EMIOENET1TXRVALID;
    input EMIOENET2DMATXSTATUSTOG;
    input EMIOENET2EXTINTIN;
    input EMIOENET2GMIICOL;
    input EMIOENET2GMIICRS;
    input EMIOENET2GMIIRXCLK;
    input [7:0] EMIOENET2GMIIRXD;
    input EMIOENET2GMIIRXDV;
    input EMIOENET2GMIIRXER;
    input EMIOENET2GMIITXCLK;
    input EMIOENET2MDIOI;
    input EMIOENET2RXWOVERFLOW;
    input EMIOENET2TXRCONTROL;
    input [7:0] EMIOENET2TXRDATA;
    input EMIOENET2TXRDATARDY;
    input EMIOENET2TXREOP;
    input EMIOENET2TXRERR;
    input EMIOENET2TXRFLUSHED;
    input EMIOENET2TXRSOP;
    input EMIOENET2TXRUNDERFLOW;
    input EMIOENET2TXRVALID;
    input EMIOENET3DMATXSTATUSTOG;
    input EMIOENET3EXTINTIN;
    input EMIOENET3GMIICOL;
    input EMIOENET3GMIICRS;
    input EMIOENET3GMIIRXCLK;
    input [7:0] EMIOENET3GMIIRXD;
    input EMIOENET3GMIIRXDV;
    input EMIOENET3GMIIRXER;
    input EMIOENET3GMIITXCLK;
    input EMIOENET3MDIOI;
    input EMIOENET3RXWOVERFLOW;
    input EMIOENET3TXRCONTROL;
    input [7:0] EMIOENET3TXRDATA;
    input EMIOENET3TXRDATARDY;
    input EMIOENET3TXREOP;
    input EMIOENET3TXRERR;
    input EMIOENET3TXRFLUSHED;
    input EMIOENET3TXRSOP;
    input EMIOENET3TXRUNDERFLOW;
    input EMIOENET3TXRVALID;
    input EMIOENETTSUCLK;
    input [1:0] EMIOGEM0TSUINCCTRL;
    input [1:0] EMIOGEM1TSUINCCTRL;
    input [1:0] EMIOGEM2TSUINCCTRL;
    input [1:0] EMIOGEM3TSUINCCTRL;
    input [95:0] EMIOGPIOI;
    input EMIOHUBPORTOVERCRNTUSB20;
    input EMIOHUBPORTOVERCRNTUSB21;
    input EMIOHUBPORTOVERCRNTUSB30;
    input EMIOHUBPORTOVERCRNTUSB31;
    input EMIOI2C0SCLI;
    input EMIOI2C0SDAI;
    input EMIOI2C1SCLI;
    input EMIOI2C1SDAI;
    input EMIOSDIO0CDN;
    input EMIOSDIO0CMDIN;
    input [7:0] EMIOSDIO0DATAIN;
    input EMIOSDIO0FBCLKIN;
    input EMIOSDIO0WP;
    input EMIOSDIO1CDN;
    input EMIOSDIO1CMDIN;
    input [7:0] EMIOSDIO1DATAIN;
    input EMIOSDIO1FBCLKIN;
    input EMIOSDIO1WP;
    input EMIOSPI0MI;
    input EMIOSPI0SCLKI;
    input EMIOSPI0SI;
    input EMIOSPI0SSIN;
    input EMIOSPI1MI;
    input EMIOSPI1SCLKI;
    input EMIOSPI1SI;
    input EMIOSPI1SSIN;
    input [2:0] EMIOTTC0CLKI;
    input [2:0] EMIOTTC1CLKI;
    input [2:0] EMIOTTC2CLKI;
    input [2:0] EMIOTTC3CLKI;
    input EMIOUART0CTSN;
    input EMIOUART0DCDN;
    input EMIOUART0DSRN;
    input EMIOUART0RIN;
    input EMIOUART0RX;
    input EMIOUART1CTSN;
    input EMIOUART1DCDN;
    input EMIOUART1DSRN;
    input EMIOUART1RIN;
    input EMIOUART1RX;
    input EMIOWDT0CLKI;
    input EMIOWDT1CLKI;
    input FMIOGEM0FIFORXCLKFROMPL;
    input FMIOGEM0FIFOTXCLKFROMPL;
    input FMIOGEM0SIGNALDETECT;
    input FMIOGEM1FIFORXCLKFROMPL;
    input FMIOGEM1FIFOTXCLKFROMPL;
    input FMIOGEM1SIGNALDETECT;
    input FMIOGEM2FIFORXCLKFROMPL;
    input FMIOGEM2FIFOTXCLKFROMPL;
    input FMIOGEM2SIGNALDETECT;
    input FMIOGEM3FIFORXCLKFROMPL;
    input FMIOGEM3FIFOTXCLKFROMPL;
    input FMIOGEM3SIGNALDETECT;
    input FMIOGEMTSUCLKFROMPL;
    input [31:0] FTMGPI;
    input [7:0] GDMAFCICLK;
    input MAXIGP0ACLK;
    input MAXIGP0ARREADY;
    input MAXIGP0AWREADY;
    input [15:0] MAXIGP0BID;
    input [1:0] MAXIGP0BRESP;
    input MAXIGP0BVALID;
    input [127:0] MAXIGP0RDATA;
    input [15:0] MAXIGP0RID;
    input MAXIGP0RLAST;
    input [1:0] MAXIGP0RRESP;
    input MAXIGP0RVALID;
    input MAXIGP0WREADY;
    input MAXIGP1ACLK;
    input MAXIGP1ARREADY;
    input MAXIGP1AWREADY;
    input [15:0] MAXIGP1BID;
    input [1:0] MAXIGP1BRESP;
    input MAXIGP1BVALID;
    input [127:0] MAXIGP1RDATA;
    input [15:0] MAXIGP1RID;
    input MAXIGP1RLAST;
    input [1:0] MAXIGP1RRESP;
    input MAXIGP1RVALID;
    input MAXIGP1WREADY;
    input MAXIGP2ACLK;
    input MAXIGP2ARREADY;
    input MAXIGP2AWREADY;
    input [15:0] MAXIGP2BID;
    input [1:0] MAXIGP2BRESP;
    input MAXIGP2BVALID;
    input [127:0] MAXIGP2RDATA;
    input [15:0] MAXIGP2RID;
    input MAXIGP2RLAST;
    input [1:0] MAXIGP2RRESP;
    input MAXIGP2RVALID;
    input MAXIGP2WREADY;
    input NFIQ0LPDRPU;
    input NFIQ1LPDRPU;
    input NIRQ0LPDRPU;
    input NIRQ1LPDRPU;
    input [7:0] PL2ADMACVLD;
    input [7:0] PL2ADMATACK;
    input [7:0] PL2GDMACVLD;
    input [7:0] PL2GDMATACK;
    input PLACECLK;
    input PLACPINACT;
    input [3:0] PLFPGASTOP;
    input [2:0] PLLAUXREFCLKFPD;
    input [1:0] PLLAUXREFCLKLPD;
    input [31:0] PLPMUGPI;
    input [3:0] PLPSAPUGICFIQ;
    input [3:0] PLPSAPUGICIRQ;
    input PLPSEVENTI;
    input [7:0] PLPSIRQ0;
    input [7:0] PLPSIRQ1;
    input PLPSTRACECLK;
    input [3:0] PLPSTRIGACK;
    input [3:0] PLPSTRIGGER;
    input [3:0] PMUERRORFROMPL;
    input PSS_ALTO_CORE_PAD_MGTRXN0IN;
    input PSS_ALTO_CORE_PAD_MGTRXN1IN;
    input PSS_ALTO_CORE_PAD_MGTRXN2IN;
    input PSS_ALTO_CORE_PAD_MGTRXN3IN;
    input PSS_ALTO_CORE_PAD_MGTRXP0IN;
    input PSS_ALTO_CORE_PAD_MGTRXP1IN;
    input PSS_ALTO_CORE_PAD_MGTRXP2IN;
    input PSS_ALTO_CORE_PAD_MGTRXP3IN;
    input PSS_ALTO_CORE_PAD_PADI;
    input PSS_ALTO_CORE_PAD_REFN0IN;
    input PSS_ALTO_CORE_PAD_REFN1IN;
    input PSS_ALTO_CORE_PAD_REFN2IN;
    input PSS_ALTO_CORE_PAD_REFN3IN;
    input PSS_ALTO_CORE_PAD_REFP0IN;
    input PSS_ALTO_CORE_PAD_REFP1IN;
    input PSS_ALTO_CORE_PAD_REFP2IN;
    input PSS_ALTO_CORE_PAD_REFP3IN;
    input RPUEVENTI0;
    input RPUEVENTI1;
    input SACEFPDACREADY;
    input [43:0] SACEFPDARADDR;
    input [1:0] SACEFPDARBAR;
    input [1:0] SACEFPDARBURST;
    input [3:0] SACEFPDARCACHE;
    input [1:0] SACEFPDARDOMAIN;
    input [5:0] SACEFPDARID;
    input [7:0] SACEFPDARLEN;
    input SACEFPDARLOCK;
    input [2:0] SACEFPDARPROT;
    input [3:0] SACEFPDARQOS;
    input [3:0] SACEFPDARREGION;
    input [2:0] SACEFPDARSIZE;
    input [3:0] SACEFPDARSNOOP;
    input [15:0] SACEFPDARUSER;
    input SACEFPDARVALID;
    input [43:0] SACEFPDAWADDR;
    input [1:0] SACEFPDAWBAR;
    input [1:0] SACEFPDAWBURST;
    input [3:0] SACEFPDAWCACHE;
    input [1:0] SACEFPDAWDOMAIN;
    input [5:0] SACEFPDAWID;
    input [7:0] SACEFPDAWLEN;
    input SACEFPDAWLOCK;
    input [2:0] SACEFPDAWPROT;
    input [3:0] SACEFPDAWQOS;
    input [3:0] SACEFPDAWREGION;
    input [2:0] SACEFPDAWSIZE;
    input [2:0] SACEFPDAWSNOOP;
    input [15:0] SACEFPDAWUSER;
    input SACEFPDAWVALID;
    input SACEFPDBREADY;
    input [127:0] SACEFPDCDDATA;
    input SACEFPDCDLAST;
    input SACEFPDCDVALID;
    input [4:0] SACEFPDCRRESP;
    input SACEFPDCRVALID;
    input SACEFPDRACK;
    input SACEFPDRREADY;
    input SACEFPDWACK;
    input [127:0] SACEFPDWDATA;
    input SACEFPDWLAST;
    input [15:0] SACEFPDWSTRB;
    input SACEFPDWUSER;
    input SACEFPDWVALID;
    input SAXIACPACLK;
    input [39:0] SAXIACPARADDR;
    input [1:0] SAXIACPARBURST;
    input [3:0] SAXIACPARCACHE;
    input [4:0] SAXIACPARID;
    input [7:0] SAXIACPARLEN;
    input SAXIACPARLOCK;
    input [2:0] SAXIACPARPROT;
    input [3:0] SAXIACPARQOS;
    input [2:0] SAXIACPARSIZE;
    input [1:0] SAXIACPARUSER;
    input SAXIACPARVALID;
    input [39:0] SAXIACPAWADDR;
    input [1:0] SAXIACPAWBURST;
    input [3:0] SAXIACPAWCACHE;
    input [4:0] SAXIACPAWID;
    input [7:0] SAXIACPAWLEN;
    input SAXIACPAWLOCK;
    input [2:0] SAXIACPAWPROT;
    input [3:0] SAXIACPAWQOS;
    input [2:0] SAXIACPAWSIZE;
    input [1:0] SAXIACPAWUSER;
    input SAXIACPAWVALID;
    input SAXIACPBREADY;
    input SAXIACPRREADY;
    input [127:0] SAXIACPWDATA;
    input SAXIACPWLAST;
    input [15:0] SAXIACPWSTRB;
    input SAXIACPWVALID;
    input [48:0] SAXIGP0ARADDR;
    input [1:0] SAXIGP0ARBURST;
    input [3:0] SAXIGP0ARCACHE;
    input [5:0] SAXIGP0ARID;
    input [7:0] SAXIGP0ARLEN;
    input SAXIGP0ARLOCK;
    input [2:0] SAXIGP0ARPROT;
    input [3:0] SAXIGP0ARQOS;
    input [2:0] SAXIGP0ARSIZE;
    input SAXIGP0ARUSER;
    input SAXIGP0ARVALID;
    input [48:0] SAXIGP0AWADDR;
    input [1:0] SAXIGP0AWBURST;
    input [3:0] SAXIGP0AWCACHE;
    input [5:0] SAXIGP0AWID;
    input [7:0] SAXIGP0AWLEN;
    input SAXIGP0AWLOCK;
    input [2:0] SAXIGP0AWPROT;
    input [3:0] SAXIGP0AWQOS;
    input [2:0] SAXIGP0AWSIZE;
    input SAXIGP0AWUSER;
    input SAXIGP0AWVALID;
    input SAXIGP0BREADY;
    input SAXIGP0RCLK;
    input SAXIGP0RREADY;
    input SAXIGP0WCLK;
    input [127:0] SAXIGP0WDATA;
    input SAXIGP0WLAST;
    input [15:0] SAXIGP0WSTRB;
    input SAXIGP0WVALID;
    input [48:0] SAXIGP1ARADDR;
    input [1:0] SAXIGP1ARBURST;
    input [3:0] SAXIGP1ARCACHE;
    input [5:0] SAXIGP1ARID;
    input [7:0] SAXIGP1ARLEN;
    input SAXIGP1ARLOCK;
    input [2:0] SAXIGP1ARPROT;
    input [3:0] SAXIGP1ARQOS;
    input [2:0] SAXIGP1ARSIZE;
    input SAXIGP1ARUSER;
    input SAXIGP1ARVALID;
    input [48:0] SAXIGP1AWADDR;
    input [1:0] SAXIGP1AWBURST;
    input [3:0] SAXIGP1AWCACHE;
    input [5:0] SAXIGP1AWID;
    input [7:0] SAXIGP1AWLEN;
    input SAXIGP1AWLOCK;
    input [2:0] SAXIGP1AWPROT;
    input [3:0] SAXIGP1AWQOS;
    input [2:0] SAXIGP1AWSIZE;
    input SAXIGP1AWUSER;
    input SAXIGP1AWVALID;
    input SAXIGP1BREADY;
    input SAXIGP1RCLK;
    input SAXIGP1RREADY;
    input SAXIGP1WCLK;
    input [127:0] SAXIGP1WDATA;
    input SAXIGP1WLAST;
    input [15:0] SAXIGP1WSTRB;
    input SAXIGP1WVALID;
    input [48:0] SAXIGP2ARADDR;
    input [1:0] SAXIGP2ARBURST;
    input [3:0] SAXIGP2ARCACHE;
    input [5:0] SAXIGP2ARID;
    input [7:0] SAXIGP2ARLEN;
    input SAXIGP2ARLOCK;
    input [2:0] SAXIGP2ARPROT;
    input [3:0] SAXIGP2ARQOS;
    input [2:0] SAXIGP2ARSIZE;
    input SAXIGP2ARUSER;
    input SAXIGP2ARVALID;
    input [48:0] SAXIGP2AWADDR;
    input [1:0] SAXIGP2AWBURST;
    input [3:0] SAXIGP2AWCACHE;
    input [5:0] SAXIGP2AWID;
    input [7:0] SAXIGP2AWLEN;
    input SAXIGP2AWLOCK;
    input [2:0] SAXIGP2AWPROT;
    input [3:0] SAXIGP2AWQOS;
    input [2:0] SAXIGP2AWSIZE;
    input SAXIGP2AWUSER;
    input SAXIGP2AWVALID;
    input SAXIGP2BREADY;
    input SAXIGP2RCLK;
    input SAXIGP2RREADY;
    input SAXIGP2WCLK;
    input [127:0] SAXIGP2WDATA;
    input SAXIGP2WLAST;
    input [15:0] SAXIGP2WSTRB;
    input SAXIGP2WVALID;
    input [48:0] SAXIGP3ARADDR;
    input [1:0] SAXIGP3ARBURST;
    input [3:0] SAXIGP3ARCACHE;
    input [5:0] SAXIGP3ARID;
    input [7:0] SAXIGP3ARLEN;
    input SAXIGP3ARLOCK;
    input [2:0] SAXIGP3ARPROT;
    input [3:0] SAXIGP3ARQOS;
    input [2:0] SAXIGP3ARSIZE;
    input SAXIGP3ARUSER;
    input SAXIGP3ARVALID;
    input [48:0] SAXIGP3AWADDR;
    input [1:0] SAXIGP3AWBURST;
    input [3:0] SAXIGP3AWCACHE;
    input [5:0] SAXIGP3AWID;
    input [7:0] SAXIGP3AWLEN;
    input SAXIGP3AWLOCK;
    input [2:0] SAXIGP3AWPROT;
    input [3:0] SAXIGP3AWQOS;
    input [2:0] SAXIGP3AWSIZE;
    input SAXIGP3AWUSER;
    input SAXIGP3AWVALID;
    input SAXIGP3BREADY;
    input SAXIGP3RCLK;
    input SAXIGP3RREADY;
    input SAXIGP3WCLK;
    input [127:0] SAXIGP3WDATA;
    input SAXIGP3WLAST;
    input [15:0] SAXIGP3WSTRB;
    input SAXIGP3WVALID;
    input [48:0] SAXIGP4ARADDR;
    input [1:0] SAXIGP4ARBURST;
    input [3:0] SAXIGP4ARCACHE;
    input [5:0] SAXIGP4ARID;
    input [7:0] SAXIGP4ARLEN;
    input SAXIGP4ARLOCK;
    input [2:0] SAXIGP4ARPROT;
    input [3:0] SAXIGP4ARQOS;
    input [2:0] SAXIGP4ARSIZE;
    input SAXIGP4ARUSER;
    input SAXIGP4ARVALID;
    input [48:0] SAXIGP4AWADDR;
    input [1:0] SAXIGP4AWBURST;
    input [3:0] SAXIGP4AWCACHE;
    input [5:0] SAXIGP4AWID;
    input [7:0] SAXIGP4AWLEN;
    input SAXIGP4AWLOCK;
    input [2:0] SAXIGP4AWPROT;
    input [3:0] SAXIGP4AWQOS;
    input [2:0] SAXIGP4AWSIZE;
    input SAXIGP4AWUSER;
    input SAXIGP4AWVALID;
    input SAXIGP4BREADY;
    input SAXIGP4RCLK;
    input SAXIGP4RREADY;
    input SAXIGP4WCLK;
    input [127:0] SAXIGP4WDATA;
    input SAXIGP4WLAST;
    input [15:0] SAXIGP4WSTRB;
    input SAXIGP4WVALID;
    input [48:0] SAXIGP5ARADDR;
    input [1:0] SAXIGP5ARBURST;
    input [3:0] SAXIGP5ARCACHE;
    input [5:0] SAXIGP5ARID;
    input [7:0] SAXIGP5ARLEN;
    input SAXIGP5ARLOCK;
    input [2:0] SAXIGP5ARPROT;
    input [3:0] SAXIGP5ARQOS;
    input [2:0] SAXIGP5ARSIZE;
    input SAXIGP5ARUSER;
    input SAXIGP5ARVALID;
    input [48:0] SAXIGP5AWADDR;
    input [1:0] SAXIGP5AWBURST;
    input [3:0] SAXIGP5AWCACHE;
    input [5:0] SAXIGP5AWID;
    input [7:0] SAXIGP5AWLEN;
    input SAXIGP5AWLOCK;
    input [2:0] SAXIGP5AWPROT;
    input [3:0] SAXIGP5AWQOS;
    input [2:0] SAXIGP5AWSIZE;
    input SAXIGP5AWUSER;
    input SAXIGP5AWVALID;
    input SAXIGP5BREADY;
    input SAXIGP5RCLK;
    input SAXIGP5RREADY;
    input SAXIGP5WCLK;
    input [127:0] SAXIGP5WDATA;
    input SAXIGP5WLAST;
    input [15:0] SAXIGP5WSTRB;
    input SAXIGP5WVALID;
    input [48:0] SAXIGP6ARADDR;
    input [1:0] SAXIGP6ARBURST;
    input [3:0] SAXIGP6ARCACHE;
    input [5:0] SAXIGP6ARID;
    input [7:0] SAXIGP6ARLEN;
    input SAXIGP6ARLOCK;
    input [2:0] SAXIGP6ARPROT;
    input [3:0] SAXIGP6ARQOS;
    input [2:0] SAXIGP6ARSIZE;
    input SAXIGP6ARUSER;
    input SAXIGP6ARVALID;
    input [48:0] SAXIGP6AWADDR;
    input [1:0] SAXIGP6AWBURST;
    input [3:0] SAXIGP6AWCACHE;
    input [5:0] SAXIGP6AWID;
    input [7:0] SAXIGP6AWLEN;
    input SAXIGP6AWLOCK;
    input [2:0] SAXIGP6AWPROT;
    input [3:0] SAXIGP6AWQOS;
    input [2:0] SAXIGP6AWSIZE;
    input SAXIGP6AWUSER;
    input SAXIGP6AWVALID;
    input SAXIGP6BREADY;
    input SAXIGP6RCLK;
    input SAXIGP6RREADY;
    input SAXIGP6WCLK;
    input [127:0] SAXIGP6WDATA;
    input SAXIGP6WLAST;
    input [15:0] SAXIGP6WSTRB;
    input SAXIGP6WVALID;
    input [59:0] STMEVENT;
endmodule

