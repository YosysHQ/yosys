// Created by cells_xtra.py from Xilinx models

module RAMB16_S1 (...);
    parameter [0:0] INIT = 1'h0;
    parameter [0:0] SRVAL = 1'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DO;
    input [13:0] ADDR;
    input [0:0] DI;
    input EN;
    (* clkbuf_sink *)
    input CLK;
    input WE;
    input SSR;
endmodule

module RAMB16_S2 (...);
    parameter [1:0] INIT = 2'h0;
    parameter [1:0] SRVAL = 2'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [1:0] DO;
    input [12:0] ADDR;
    input [1:0] DI;
    input EN;
    (* clkbuf_sink *)
    input CLK;
    input WE;
    input SSR;
endmodule

module RAMB16_S4 (...);
    parameter [3:0] INIT = 4'h0;
    parameter [3:0] SRVAL = 4'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [3:0] DO;
    input [11:0] ADDR;
    input [3:0] DI;
    input EN;
    (* clkbuf_sink *)
    input CLK;
    input WE;
    input SSR;
endmodule

module RAMB16_S9 (...);
    parameter [8:0] INIT = 9'h0;
    parameter [8:0] SRVAL = 9'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [7:0] DO;
    output [0:0] DOP;
    input [10:0] ADDR;
    input [7:0] DI;
    input [0:0] DIP;
    input EN;
    (* clkbuf_sink *)
    input CLK;
    input WE;
    input SSR;
endmodule

module RAMB16_S18 (...);
    parameter [17:0] INIT = 18'h0;
    parameter [17:0] SRVAL = 18'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [15:0] DO;
    output [1:0] DOP;
    input [9:0] ADDR;
    input [15:0] DI;
    input [1:0] DIP;
    input EN;
    (* clkbuf_sink *)
    input CLK;
    input WE;
    input SSR;
endmodule

module RAMB16_S36 (...);
    parameter [35:0] INIT = 36'h0;
    parameter [35:0] SRVAL = 36'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [31:0] DO;
    output [3:0] DOP;
    input [8:0] ADDR;
    input [31:0] DI;
    input [3:0] DIP;
    input EN;
    (* clkbuf_sink *)
    input CLK;
    input WE;
    input SSR;
endmodule

module RAMB16_S1_S1 (...);
    parameter [0:0] INIT_A = 1'h0;
    parameter [0:0] INIT_B = 1'h0;
    parameter [0:0] SRVAL_A = 1'h0;
    parameter [0:0] SRVAL_B = 1'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DOA;
    input [13:0] ADDRA;
    input [0:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [0:0] DOB;
    input [13:0] ADDRB;
    input [0:0] DIB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S1_S2 (...);
    parameter [0:0] INIT_A = 1'h0;
    parameter [1:0] INIT_B = 2'h0;
    parameter [0:0] SRVAL_A = 1'h0;
    parameter [1:0] SRVAL_B = 2'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DOA;
    input [13:0] ADDRA;
    input [0:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [1:0] DOB;
    input [12:0] ADDRB;
    input [1:0] DIB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S1_S4 (...);
    parameter [0:0] INIT_A = 1'h0;
    parameter [3:0] INIT_B = 4'h0;
    parameter [0:0] SRVAL_A = 1'h0;
    parameter [3:0] SRVAL_B = 4'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DOA;
    input [13:0] ADDRA;
    input [0:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [3:0] DOB;
    input [11:0] ADDRB;
    input [3:0] DIB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S1_S9 (...);
    parameter [0:0] INIT_A = 1'h0;
    parameter [8:0] INIT_B = 9'h0;
    parameter [0:0] SRVAL_A = 1'h0;
    parameter [8:0] SRVAL_B = 9'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DOA;
    input [13:0] ADDRA;
    input [0:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [7:0] DOB;
    output [0:0] DOPB;
    input [10:0] ADDRB;
    input [7:0] DIB;
    input [0:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S1_S18 (...);
    parameter [0:0] INIT_A = 1'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter [0:0] SRVAL_A = 1'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DOA;
    input [13:0] ADDRA;
    input [0:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [15:0] DOB;
    output [1:0] DOPB;
    input [9:0] ADDRB;
    input [15:0] DIB;
    input [1:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S1_S36 (...);
    parameter [0:0] INIT_A = 1'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter [0:0] SRVAL_A = 1'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [0:0] DOA;
    input [13:0] ADDRA;
    input [0:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [31:0] DOB;
    output [3:0] DOPB;
    input [8:0] ADDRB;
    input [31:0] DIB;
    input [3:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S2_S2 (...);
    parameter [1:0] INIT_A = 2'h0;
    parameter [1:0] INIT_B = 2'h0;
    parameter [1:0] SRVAL_A = 2'h0;
    parameter [1:0] SRVAL_B = 2'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [1:0] DOA;
    input [12:0] ADDRA;
    input [1:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [1:0] DOB;
    input [12:0] ADDRB;
    input [1:0] DIB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S2_S4 (...);
    parameter [1:0] INIT_A = 2'h0;
    parameter [3:0] INIT_B = 4'h0;
    parameter [1:0] SRVAL_A = 2'h0;
    parameter [3:0] SRVAL_B = 4'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [1:0] DOA;
    input [12:0] ADDRA;
    input [1:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [3:0] DOB;
    input [11:0] ADDRB;
    input [3:0] DIB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S2_S9 (...);
    parameter [1:0] INIT_A = 2'h0;
    parameter [8:0] INIT_B = 9'h0;
    parameter [1:0] SRVAL_A = 2'h0;
    parameter [8:0] SRVAL_B = 9'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [1:0] DOA;
    input [12:0] ADDRA;
    input [1:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [7:0] DOB;
    output [0:0] DOPB;
    input [10:0] ADDRB;
    input [7:0] DIB;
    input [0:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S2_S18 (...);
    parameter [1:0] INIT_A = 2'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter [1:0] SRVAL_A = 2'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [1:0] DOA;
    input [12:0] ADDRA;
    input [1:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [15:0] DOB;
    output [1:0] DOPB;
    input [9:0] ADDRB;
    input [15:0] DIB;
    input [1:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S2_S36 (...);
    parameter [1:0] INIT_A = 2'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter [1:0] SRVAL_A = 2'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [1:0] DOA;
    input [12:0] ADDRA;
    input [1:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [31:0] DOB;
    output [3:0] DOPB;
    input [8:0] ADDRB;
    input [31:0] DIB;
    input [3:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S4_S4 (...);
    parameter [3:0] INIT_A = 4'h0;
    parameter [3:0] INIT_B = 4'h0;
    parameter [3:0] SRVAL_A = 4'h0;
    parameter [3:0] SRVAL_B = 4'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [3:0] DOA;
    input [11:0] ADDRA;
    input [3:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [3:0] DOB;
    input [11:0] ADDRB;
    input [3:0] DIB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S4_S9 (...);
    parameter [3:0] INIT_A = 4'h0;
    parameter [8:0] INIT_B = 9'h0;
    parameter [3:0] SRVAL_A = 4'h0;
    parameter [8:0] SRVAL_B = 9'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [3:0] DOA;
    input [11:0] ADDRA;
    input [3:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [7:0] DOB;
    output [0:0] DOPB;
    input [10:0] ADDRB;
    input [7:0] DIB;
    input [0:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S4_S18 (...);
    parameter [3:0] INIT_A = 4'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter [3:0] SRVAL_A = 4'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [3:0] DOA;
    input [11:0] ADDRA;
    input [3:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [15:0] DOB;
    output [1:0] DOPB;
    input [9:0] ADDRB;
    input [15:0] DIB;
    input [1:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S4_S36 (...);
    parameter [3:0] INIT_A = 4'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter [3:0] SRVAL_A = 4'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [3:0] DOA;
    input [11:0] ADDRA;
    input [3:0] DIA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [31:0] DOB;
    output [3:0] DOPB;
    input [8:0] ADDRB;
    input [31:0] DIB;
    input [3:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S9_S9 (...);
    parameter [8:0] INIT_A = 9'h0;
    parameter [8:0] INIT_B = 9'h0;
    parameter [8:0] SRVAL_A = 9'h0;
    parameter [8:0] SRVAL_B = 9'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [7:0] DOA;
    output [0:0] DOPA;
    input [10:0] ADDRA;
    input [7:0] DIA;
    input [0:0] DIPA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [7:0] DOB;
    output [0:0] DOPB;
    input [10:0] ADDRB;
    input [7:0] DIB;
    input [0:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S9_S18 (...);
    parameter [8:0] INIT_A = 9'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter [8:0] SRVAL_A = 9'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [7:0] DOA;
    output [0:0] DOPA;
    input [10:0] ADDRA;
    input [7:0] DIA;
    input [0:0] DIPA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [15:0] DOB;
    output [1:0] DOPB;
    input [9:0] ADDRB;
    input [15:0] DIB;
    input [1:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S9_S36 (...);
    parameter [8:0] INIT_A = 9'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter [8:0] SRVAL_A = 9'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [7:0] DOA;
    output [0:0] DOPA;
    input [10:0] ADDRA;
    input [7:0] DIA;
    input [0:0] DIPA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [31:0] DOB;
    output [3:0] DOPB;
    input [8:0] ADDRB;
    input [31:0] DIB;
    input [3:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S18_S18 (...);
    parameter [17:0] INIT_A = 18'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter [17:0] SRVAL_A = 18'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [15:0] DOA;
    output [1:0] DOPA;
    input [9:0] ADDRA;
    input [15:0] DIA;
    input [1:0] DIPA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [15:0] DOB;
    output [1:0] DOPB;
    input [9:0] ADDRB;
    input [15:0] DIB;
    input [1:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S18_S36 (...);
    parameter [17:0] INIT_A = 18'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter [17:0] SRVAL_A = 18'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [15:0] DOA;
    output [1:0] DOPA;
    input [9:0] ADDRA;
    input [15:0] DIA;
    input [1:0] DIPA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [31:0] DOB;
    output [3:0] DOPB;
    input [8:0] ADDRB;
    input [31:0] DIB;
    input [3:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16_S36_S36 (...);
    parameter [35:0] INIT_A = 36'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output [31:0] DOA;
    output [3:0] DOPA;
    input [8:0] ADDRA;
    input [31:0] DIA;
    input [3:0] DIPA;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input WEA;
    input SSRA;
    output [31:0] DOB;
    output [3:0] DOPB;
    input [8:0] ADDRB;
    input [31:0] DIB;
    input [3:0] DIPB;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input WEB;
    input SSRB;
endmodule

module RAMB16BWE_S18 (...);
    parameter [17:0] INIT = 18'h0;
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [17:0] SRVAL = 18'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    output [15:0] DO;
    output [1:0] DOP;
    (* clkbuf_sink *)
    input CLK;
    input EN;
    input SSR;
    input [1:0] WE;
    input [15:0] DI;
    input [1:0] DIP;
    input [9:0] ADDR;
endmodule

module RAMB16BWE_S36 (...);
    parameter [35:0] INIT = 36'h0;
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [35:0] SRVAL = 36'h0;
    parameter WRITE_MODE = "WRITE_FIRST";
    output [31:0] DO;
    output [3:0] DOP;
    (* clkbuf_sink *)
    input CLK;
    input EN;
    input SSR;
    input [3:0] WE;
    input [31:0] DI;
    input [3:0] DIP;
    input [8:0] ADDR;
endmodule

module RAMB16BWE_S18_S9 (...);
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [17:0] INIT_A = 18'h0;
    parameter [8:0] INIT_B = 9'h0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [17:0] SRVAL_A = 18'h0;
    parameter [8:0] SRVAL_B = 9'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [15:0] DOA;
    output [7:0] DOB;
    output [1:0] DOPA;
    output [0:0] DOPB;
    (* clkbuf_sink *)
    input CLKA;
    (* clkbuf_sink *)
    input CLKB;
    input ENA;
    input ENB;
    input SSRA;
    input SSRB;
    input WEB;
    input [1:0] WEA;
    input [15:0] DIA;
    input [7:0] DIB;
    input [1:0] DIPA;
    input [0:0] DIPB;
    input [9:0] ADDRA;
    input [10:0] ADDRB;
endmodule

module RAMB16BWE_S18_S18 (...);
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [17:0] INIT_A = 18'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [17:0] SRVAL_A = 18'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [15:0] DOA;
    output [15:0] DOB;
    output [1:0] DOPA;
    output [1:0] DOPB;
    (* clkbuf_sink *)
    input CLKA;
    (* clkbuf_sink *)
    input CLKB;
    input ENA;
    input ENB;
    input SSRA;
    input SSRB;
    input [1:0] WEB;
    input [1:0] WEA;
    input [15:0] DIA;
    input [15:0] DIB;
    input [1:0] DIPA;
    input [1:0] DIPB;
    input [9:0] ADDRA;
    input [9:0] ADDRB;
endmodule

module RAMB16BWE_S36_S9 (...);
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [35:0] INIT_A = 36'h0;
    parameter [8:0] INIT_B = 9'h0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [8:0] SRVAL_B = 9'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [31:0] DOA;
    output [3:0] DOPA;
    output [7:0] DOB;
    output [0:0] DOPB;
    (* clkbuf_sink *)
    input CLKA;
    (* clkbuf_sink *)
    input CLKB;
    input ENA;
    input ENB;
    input SSRA;
    input SSRB;
    input [3:0] WEA;
    input WEB;
    input [31:0] DIA;
    input [3:0] DIPA;
    input [7:0] DIB;
    input [0:0] DIPB;
    input [8:0] ADDRA;
    input [10:0] ADDRB;
endmodule

module RAMB16BWE_S36_S18 (...);
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [35:0] INIT_A = 36'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [31:0] DOA;
    output [3:0] DOPA;
    output [15:0] DOB;
    output [1:0] DOPB;
    (* clkbuf_sink *)
    input CLKA;
    (* clkbuf_sink *)
    input CLKB;
    input ENA;
    input ENB;
    input SSRA;
    input SSRB;
    input [3:0] WEA;
    input [1:0] WEB;
    input [31:0] DIA;
    input [3:0] DIPA;
    input [15:0] DIB;
    input [1:0] DIPB;
    input [8:0] ADDRA;
    input [9:0] ADDRB;
endmodule

module RAMB16BWE_S36_S36 (...);
    parameter [255:0] INITP_00 = 256'h0;
    parameter [255:0] INITP_01 = 256'h0;
    parameter [255:0] INITP_02 = 256'h0;
    parameter [255:0] INITP_03 = 256'h0;
    parameter [255:0] INITP_04 = 256'h0;
    parameter [255:0] INITP_05 = 256'h0;
    parameter [255:0] INITP_06 = 256'h0;
    parameter [255:0] INITP_07 = 256'h0;
    parameter [255:0] INIT_00 = 256'h0;
    parameter [255:0] INIT_01 = 256'h0;
    parameter [255:0] INIT_02 = 256'h0;
    parameter [255:0] INIT_03 = 256'h0;
    parameter [255:0] INIT_04 = 256'h0;
    parameter [255:0] INIT_05 = 256'h0;
    parameter [255:0] INIT_06 = 256'h0;
    parameter [255:0] INIT_07 = 256'h0;
    parameter [255:0] INIT_08 = 256'h0;
    parameter [255:0] INIT_09 = 256'h0;
    parameter [255:0] INIT_0A = 256'h0;
    parameter [255:0] INIT_0B = 256'h0;
    parameter [255:0] INIT_0C = 256'h0;
    parameter [255:0] INIT_0D = 256'h0;
    parameter [255:0] INIT_0E = 256'h0;
    parameter [255:0] INIT_0F = 256'h0;
    parameter [255:0] INIT_10 = 256'h0;
    parameter [255:0] INIT_11 = 256'h0;
    parameter [255:0] INIT_12 = 256'h0;
    parameter [255:0] INIT_13 = 256'h0;
    parameter [255:0] INIT_14 = 256'h0;
    parameter [255:0] INIT_15 = 256'h0;
    parameter [255:0] INIT_16 = 256'h0;
    parameter [255:0] INIT_17 = 256'h0;
    parameter [255:0] INIT_18 = 256'h0;
    parameter [255:0] INIT_19 = 256'h0;
    parameter [255:0] INIT_1A = 256'h0;
    parameter [255:0] INIT_1B = 256'h0;
    parameter [255:0] INIT_1C = 256'h0;
    parameter [255:0] INIT_1D = 256'h0;
    parameter [255:0] INIT_1E = 256'h0;
    parameter [255:0] INIT_1F = 256'h0;
    parameter [255:0] INIT_20 = 256'h0;
    parameter [255:0] INIT_21 = 256'h0;
    parameter [255:0] INIT_22 = 256'h0;
    parameter [255:0] INIT_23 = 256'h0;
    parameter [255:0] INIT_24 = 256'h0;
    parameter [255:0] INIT_25 = 256'h0;
    parameter [255:0] INIT_26 = 256'h0;
    parameter [255:0] INIT_27 = 256'h0;
    parameter [255:0] INIT_28 = 256'h0;
    parameter [255:0] INIT_29 = 256'h0;
    parameter [255:0] INIT_2A = 256'h0;
    parameter [255:0] INIT_2B = 256'h0;
    parameter [255:0] INIT_2C = 256'h0;
    parameter [255:0] INIT_2D = 256'h0;
    parameter [255:0] INIT_2E = 256'h0;
    parameter [255:0] INIT_2F = 256'h0;
    parameter [255:0] INIT_30 = 256'h0;
    parameter [255:0] INIT_31 = 256'h0;
    parameter [255:0] INIT_32 = 256'h0;
    parameter [255:0] INIT_33 = 256'h0;
    parameter [255:0] INIT_34 = 256'h0;
    parameter [255:0] INIT_35 = 256'h0;
    parameter [255:0] INIT_36 = 256'h0;
    parameter [255:0] INIT_37 = 256'h0;
    parameter [255:0] INIT_38 = 256'h0;
    parameter [255:0] INIT_39 = 256'h0;
    parameter [255:0] INIT_3A = 256'h0;
    parameter [255:0] INIT_3B = 256'h0;
    parameter [255:0] INIT_3C = 256'h0;
    parameter [255:0] INIT_3D = 256'h0;
    parameter [255:0] INIT_3E = 256'h0;
    parameter [255:0] INIT_3F = 256'h0;
    parameter [35:0] INIT_A = 36'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [31:0] DOA;
    output [3:0] DOPA;
    output [31:0] DOB;
    output [3:0] DOPB;
    (* clkbuf_sink *)
    input CLKA;
    (* clkbuf_sink *)
    input CLKB;
    input ENA;
    input ENB;
    input SSRA;
    input SSRB;
    input [3:0] WEA;
    input [3:0] WEB;
    input [31:0] DIA;
    input [3:0] DIPA;
    input [31:0] DIB;
    input [3:0] DIPB;
    input [8:0] ADDRA;
    input [8:0] ADDRB;
endmodule

module RAMB16BWER (...);
    parameter integer DATA_WIDTH_A = 0;
    parameter integer DATA_WIDTH_B = 0;
    parameter integer DOA_REG = 0;
    parameter integer DOB_REG = 0;
    parameter EN_RSTRAM_A = "TRUE";
    parameter EN_RSTRAM_B = "TRUE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [35:0] INIT_A = 36'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter INIT_FILE = "NONE";
    parameter RSTTYPE = "SYNC";
    parameter RST_PRIORITY_A = "CE";
    parameter RST_PRIORITY_B = "CE";
    parameter SETUP_ALL = 1000;
    parameter SETUP_READ_FIRST = 3000;
    parameter SIM_DEVICE = "SPARTAN3ADSP";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [31:0] DOA;
    output [31:0] DOB;
    output [3:0] DOPA;
    output [3:0] DOPB;
    input [13:0] ADDRA;
    input [13:0] ADDRB;
    (* clkbuf_sink *)
    input CLKA;
    (* clkbuf_sink *)
    input CLKB;
    input [31:0] DIA;
    input [31:0] DIB;
    input [3:0] DIPA;
    input [3:0] DIPB;
    input ENA;
    input ENB;
    input REGCEA;
    input REGCEB;
    input RSTA;
    input RSTB;
    input [3:0] WEA;
    input [3:0] WEB;
endmodule

module RAMB8BWER (...);
    parameter integer DATA_WIDTH_A = 0;
    parameter integer DATA_WIDTH_B = 0;
    parameter integer DOA_REG = 0;
    parameter integer DOB_REG = 0;
    parameter EN_RSTRAM_A = "TRUE";
    parameter EN_RSTRAM_B = "TRUE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [17:0] INIT_A = 18'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter INIT_FILE = "NONE";
    parameter RAM_MODE = "TDP";
    parameter RSTTYPE = "SYNC";
    parameter RST_PRIORITY_A = "CE";
    parameter RST_PRIORITY_B = "CE";
    parameter SETUP_ALL = 1000;
    parameter SETUP_READ_FIRST = 3000;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [17:0] SRVAL_A = 18'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    output [15:0] DOADO;
    output [15:0] DOBDO;
    output [1:0] DOPADOP;
    output [1:0] DOPBDOP;
    input [12:0] ADDRAWRADDR;
    input [12:0] ADDRBRDADDR;
    (* clkbuf_sink *)
    input CLKAWRCLK;
    (* clkbuf_sink *)
    input CLKBRDCLK;
    input [15:0] DIADI;
    input [15:0] DIBDI;
    input [1:0] DIPADIP;
    input [1:0] DIPBDIP;
    input ENAWREN;
    input ENBRDEN;
    input REGCEA;
    input REGCEBREGCE;
    input RSTA;
    input RSTBRST;
    input [1:0] WEAWEL;
    input [1:0] WEBWEU;
endmodule

module FIFO16 (...);
    parameter [11:0] ALMOST_FULL_OFFSET = 12'h080;
    parameter [11:0] ALMOST_EMPTY_OFFSET = 12'h080;
    parameter integer DATA_WIDTH = 36;
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [31:0] DO;
    output [3:0] DOP;
    output EMPTY;
    output FULL;
    output [11:0] RDCOUNT;
    output RDERR;
    output [11:0] WRCOUNT;
    output WRERR;
    input [31:0] DI;
    input [3:0] DIP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RST;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module RAMB16 (...);
    parameter integer DOA_REG = 0;
    parameter integer DOB_REG = 0;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [35:0] INIT_A = 36'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter INIT_FILE = "NONE";
    parameter INVERT_CLK_DOA_REG = "FALSE";
    parameter INVERT_CLK_DOB_REG = "FALSE";
    parameter RAM_EXTENSION_A = "NONE";
    parameter RAM_EXTENSION_B = "NONE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output CASCADEOUTA;
    output CASCADEOUTB;
    output [31:0] DOA;
    output [31:0] DOB;
    output [3:0] DOPA;
    output [3:0] DOPB;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input SSRA;
    input CASCADEINA;
    input REGCEA;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input SSRB;
    input CASCADEINB;
    input REGCEB;
    input [14:0] ADDRA;
    input [14:0] ADDRB;
    input [31:0] DIA;
    input [31:0] DIB;
    input [3:0] DIPA;
    input [3:0] DIPB;
    input [3:0] WEA;
    input [3:0] WEB;
endmodule

module RAMB32_S64_ECC (...);
    parameter DO_REG = 0;
    parameter SIM_COLLISION_CHECK = "ALL";
    output [1:0] STATUS;
    output [63:0] DO;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input SSR;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [63:0] DI;
    input [8:0] RDADDR;
    input [8:0] WRADDR;
endmodule

module FIFO18 (...);
    parameter [11:0] ALMOST_EMPTY_OFFSET = 12'h080;
    parameter [11:0] ALMOST_FULL_OFFSET = 12'h080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_SYN = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter SIM_MODE = "SAFE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [15:0] DO;
    output [1:0] DOP;
    output EMPTY;
    output FULL;
    output [11:0] RDCOUNT;
    output RDERR;
    output [11:0] WRCOUNT;
    output WRERR;
    input [15:0] DI;
    input [1:0] DIP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RST;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module FIFO18_36 (...);
    parameter [8:0] ALMOST_EMPTY_OFFSET = 9'h080;
    parameter [8:0] ALMOST_FULL_OFFSET = 9'h080;
    parameter integer DO_REG = 1;
    parameter EN_SYN = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter SIM_MODE = "SAFE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [31:0] DO;
    output [3:0] DOP;
    output EMPTY;
    output FULL;
    output [8:0] RDCOUNT;
    output RDERR;
    output [8:0] WRCOUNT;
    output WRERR;
    input [31:0] DI;
    input [3:0] DIP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RST;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module FIFO36 (...);
    parameter [12:0] ALMOST_EMPTY_OFFSET = 13'h080;
    parameter [12:0] ALMOST_FULL_OFFSET = 13'h080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_SYN = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter SIM_MODE = "SAFE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [31:0] DO;
    output [3:0] DOP;
    output EMPTY;
    output FULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output [12:0] WRCOUNT;
    output WRERR;
    input [31:0] DI;
    input [3:0] DIP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RST;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module FIFO36_72 (...);
    parameter [8:0] ALMOST_EMPTY_OFFSET = 9'h080;
    parameter [8:0] ALMOST_FULL_OFFSET = 9'h080;
    parameter integer DO_REG = 1;
    parameter EN_ECC_WRITE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_SYN = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter SIM_MODE = "SAFE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output DBITERR;
    output [63:0] DO;
    output [7:0] DOP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output [8:0] RDCOUNT;
    output RDERR;
    output SBITERR;
    output [8:0] WRCOUNT;
    output WRERR;
    input [63:0] DI;
    input [7:0] DIP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RST;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module RAMB18 (...);
    parameter integer DOA_REG = 0;
    parameter integer DOB_REG = 0;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [17:0] INIT_A = 18'h0;
    parameter [17:0] INIT_B = 18'h0;
    parameter INIT_FILE = "NONE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SIM_MODE = "SAFE";
    parameter [17:0] SRVAL_A = 18'h0;
    parameter [17:0] SRVAL_B = 18'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [15:0] DOA;
    output [15:0] DOB;
    output [1:0] DOPA;
    output [1:0] DOPB;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input SSRA;
    input REGCEA;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input SSRB;
    input REGCEB;
    input [13:0] ADDRA;
    input [13:0] ADDRB;
    input [15:0] DIA;
    input [15:0] DIB;
    input [1:0] DIPA;
    input [1:0] DIPB;
    input [1:0] WEA;
    input [1:0] WEB;
endmodule

module RAMB36 (...);
    parameter integer DOA_REG = 0;
    parameter integer DOB_REG = 0;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [35:0] INIT_A = 36'h0;
    parameter [35:0] INIT_B = 36'h0;
    parameter INIT_FILE = "NONE";
    parameter RAM_EXTENSION_A = "NONE";
    parameter RAM_EXTENSION_B = "NONE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SIM_MODE = "SAFE";
    parameter [35:0] SRVAL_A = 36'h0;
    parameter [35:0] SRVAL_B = 36'h0;
    parameter WRITE_MODE_A = "WRITE_FIRST";
    parameter WRITE_MODE_B = "WRITE_FIRST";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output CASCADEOUTLATA;
    output CASCADEOUTREGA;
    output CASCADEOUTLATB;
    output CASCADEOUTREGB;
    output [31:0] DOA;
    output [31:0] DOB;
    output [3:0] DOPA;
    output [3:0] DOPB;
    input ENA;
    (* clkbuf_sink *)
    input CLKA;
    input SSRA;
    input CASCADEINLATA;
    input CASCADEINREGA;
    input REGCEA;
    input ENB;
    (* clkbuf_sink *)
    input CLKB;
    input SSRB;
    input CASCADEINLATB;
    input CASCADEINREGB;
    input REGCEB;
    input [15:0] ADDRA;
    input [15:0] ADDRB;
    input [31:0] DIA;
    input [31:0] DIB;
    input [3:0] DIPA;
    input [3:0] DIPB;
    input [3:0] WEA;
    input [3:0] WEB;
endmodule

module RAMB18SDP (...);
    parameter integer DO_REG = 0;
    parameter [35:0] INIT = 36'h0;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_FILE = "NONE";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SIM_MODE = "SAFE";
    parameter [35:0] SRVAL = 36'h0;
    output [31:0] DO;
    output [3:0] DOP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input REGCE;
    input SSR;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [8:0] WRADDR;
    input [8:0] RDADDR;
    input [31:0] DI;
    input [3:0] DIP;
    input [3:0] WE;
endmodule

module RAMB36SDP (...);
    parameter integer DO_REG = 0;
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_SCRUB = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter [71:0] INIT = 72'h0;
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_FILE = "NONE";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SIM_MODE = "SAFE";
    parameter [71:0] SRVAL = 72'h0;
    output DBITERR;
    output SBITERR;
    output [63:0] DO;
    output [7:0] DOP;
    output [7:0] ECCPARITY;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input REGCE;
    input SSR;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [8:0] WRADDR;
    input [8:0] RDADDR;
    input [63:0] DI;
    input [7:0] DIP;
    input [7:0] WE;
endmodule

module FIFO18E1 (...);
    parameter ALMOST_EMPTY_OFFSET = 13'h0080;
    parameter ALMOST_FULL_OFFSET = 13'h0080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_SYN = "FALSE";
    parameter FIFO_MODE = "FIFO18";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter INIT = 36'h0;
    parameter SIM_DEVICE = "VIRTEX6";
    parameter SRVAL = 36'h0;
    parameter IS_RDCLK_INVERTED = 1'b0;
    parameter IS_RDEN_INVERTED = 1'b0;
    parameter IS_RSTREG_INVERTED = 1'b0;
    parameter IS_RST_INVERTED = 1'b0;
    parameter IS_WRCLK_INVERTED = 1'b0;
    parameter IS_WREN_INVERTED = 1'b0;
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [31:0] DO;
    output [3:0] DOP;
    output EMPTY;
    output FULL;
    output [11:0] RDCOUNT;
    output RDERR;
    output [11:0] WRCOUNT;
    output WRERR;
    input [31:0] DI;
    input [3:0] DIP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module FIFO36E1 (...);
    parameter ALMOST_EMPTY_OFFSET = 13'h0080;
    parameter ALMOST_FULL_OFFSET = 13'h0080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter EN_SYN = "FALSE";
    parameter FIFO_MODE = "FIFO36";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter INIT = 72'h0;
    parameter SIM_DEVICE = "VIRTEX6";
    parameter SRVAL = 72'h0;
    parameter IS_RDCLK_INVERTED = 1'b0;
    parameter IS_RDEN_INVERTED = 1'b0;
    parameter IS_RSTREG_INVERTED = 1'b0;
    parameter IS_RST_INVERTED = 1'b0;
    parameter IS_WRCLK_INVERTED = 1'b0;
    parameter IS_WREN_INVERTED = 1'b0;
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output DBITERR;
    output [63:0] DO;
    output [7:0] DOP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output SBITERR;
    output [12:0] WRCOUNT;
    output WRERR;
    input [63:0] DI;
    input [7:0] DIP;
    input INJECTDBITERR;
    input INJECTSBITERR;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module FIFO18E2 (...);
    parameter CASCADE_ORDER = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter [35:0] INIT = 36'h000000000;
    parameter [0:0] IS_RDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RDEN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_WRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_WREN_INVERTED = 1'b0;
    parameter integer PROG_EMPTY_THRESH = 256;
    parameter integer PROG_FULL_THRESH = 256;
    parameter RDCOUNT_TYPE = "RAW_PNTR";
    parameter integer READ_WIDTH = 4;
    parameter REGISTER_MODE = "UNREGISTERED";
    parameter RSTREG_PRIORITY = "RSTREG";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [35:0] SRVAL = 36'h000000000;
    parameter WRCOUNT_TYPE = "RAW_PNTR";
    parameter integer WRITE_WIDTH = 4;
    output [31:0] CASDOUT;
    output [3:0] CASDOUTP;
    output CASNXTEMPTY;
    output CASPRVRDEN;
    output [31:0] DOUT;
    output [3:0] DOUTP;
    output EMPTY;
    output FULL;
    output PROGEMPTY;
    output PROGFULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output RDRSTBUSY;
    output [12:0] WRCOUNT;
    output WRERR;
    output WRRSTBUSY;
    input [31:0] CASDIN;
    input [3:0] CASDINP;
    input CASDOMUX;
    input CASDOMUXEN;
    input CASNXTRDEN;
    input CASOREGIMUX;
    input CASOREGIMUXEN;
    input CASPRVEMPTY;
    input [31:0] DIN;
    input [3:0] DINP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    input SLEEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module FIFO36E2 (...);
    parameter CASCADE_ORDER = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter EN_ECC_PIPE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter [71:0] INIT = 72'h000000000000000000;
    parameter [0:0] IS_RDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RDEN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_WRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_WREN_INVERTED = 1'b0;
    parameter integer PROG_EMPTY_THRESH = 256;
    parameter integer PROG_FULL_THRESH = 256;
    parameter RDCOUNT_TYPE = "RAW_PNTR";
    parameter integer READ_WIDTH = 4;
    parameter REGISTER_MODE = "UNREGISTERED";
    parameter RSTREG_PRIORITY = "RSTREG";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [71:0] SRVAL = 72'h000000000000000000;
    parameter WRCOUNT_TYPE = "RAW_PNTR";
    parameter integer WRITE_WIDTH = 4;
    output [63:0] CASDOUT;
    output [7:0] CASDOUTP;
    output CASNXTEMPTY;
    output CASPRVRDEN;
    output DBITERR;
    output [63:0] DOUT;
    output [7:0] DOUTP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output PROGEMPTY;
    output PROGFULL;
    output [13:0] RDCOUNT;
    output RDERR;
    output RDRSTBUSY;
    output SBITERR;
    output [13:0] WRCOUNT;
    output WRERR;
    output WRRSTBUSY;
    input [63:0] CASDIN;
    input [7:0] CASDINP;
    input CASDOMUX;
    input CASDOMUXEN;
    input CASNXTRDEN;
    input CASOREGIMUX;
    input CASOREGIMUXEN;
    input CASPRVEMPTY;
    input [63:0] DIN;
    input [7:0] DINP;
    input INJECTDBITERR;
    input INJECTSBITERR;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    input SLEEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module RAMB18E2 (...);
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter integer DOA_REG = 1;
    parameter integer DOB_REG = 1;
    parameter ENADDRENA = "FALSE";
    parameter ENADDRENB = "FALSE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [17:0] INIT_A = 18'h00000;
    parameter [17:0] INIT_B = 18'h00000;
    parameter INIT_FILE = "NONE";
    parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
    parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
    parameter RDADDRCHANGEA = "FALSE";
    parameter RDADDRCHANGEB = "FALSE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter RSTREG_PRIORITY_A = "RSTREG";
    parameter RSTREG_PRIORITY_B = "RSTREG";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [17:0] SRVAL_A = 18'h00000;
    parameter [17:0] SRVAL_B = 18'h00000;
    parameter WRITE_MODE_A = "NO_CHANGE";
    parameter WRITE_MODE_B = "NO_CHANGE";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [15:0] CASDOUTA;
    output [15:0] CASDOUTB;
    output [1:0] CASDOUTPA;
    output [1:0] CASDOUTPB;
    output [15:0] DOUTADOUT;
    output [15:0] DOUTBDOUT;
    output [1:0] DOUTPADOUTP;
    output [1:0] DOUTPBDOUTP;
    input [13:0] ADDRARDADDR;
    input [13:0] ADDRBWRADDR;
    input ADDRENA;
    input ADDRENB;
    input CASDIMUXA;
    input CASDIMUXB;
    input [15:0] CASDINA;
    input [15:0] CASDINB;
    input [1:0] CASDINPA;
    input [1:0] CASDINPB;
    input CASDOMUXA;
    input CASDOMUXB;
    input CASDOMUXEN_A;
    input CASDOMUXEN_B;
    input CASOREGIMUXA;
    input CASOREGIMUXB;
    input CASOREGIMUXEN_A;
    input CASOREGIMUXEN_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKARDCLK_INVERTED" *)
    input CLKARDCLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKBWRCLK_INVERTED" *)
    input CLKBWRCLK;
    input [15:0] DINADIN;
    input [15:0] DINBDIN;
    input [1:0] DINPADINP;
    input [1:0] DINPBDINP;
    (* invertible_pin = "IS_ENARDEN_INVERTED" *)
    input ENARDEN;
    (* invertible_pin = "IS_ENBWREN_INVERTED" *)
    input ENBWREN;
    input REGCEAREGCE;
    input REGCEB;
    (* invertible_pin = "IS_RSTRAMARSTRAM_INVERTED" *)
    input RSTRAMARSTRAM;
    (* invertible_pin = "IS_RSTRAMB_INVERTED" *)
    input RSTRAMB;
    (* invertible_pin = "IS_RSTREGARSTREG_INVERTED" *)
    input RSTREGARSTREG;
    (* invertible_pin = "IS_RSTREGB_INVERTED" *)
    input RSTREGB;
    input SLEEP;
    input [1:0] WEA;
    input [3:0] WEBWE;
endmodule

module RAMB36E2 (...);
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter integer DOA_REG = 1;
    parameter integer DOB_REG = 1;
    parameter ENADDRENA = "FALSE";
    parameter ENADDRENB = "FALSE";
    parameter EN_ECC_PIPE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [35:0] INIT_A = 36'h000000000;
    parameter [35:0] INIT_B = 36'h000000000;
    parameter INIT_FILE = "NONE";
    parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
    parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
    parameter RDADDRCHANGEA = "FALSE";
    parameter RDADDRCHANGEB = "FALSE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter RSTREG_PRIORITY_A = "RSTREG";
    parameter RSTREG_PRIORITY_B = "RSTREG";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [35:0] SRVAL_A = 36'h000000000;
    parameter [35:0] SRVAL_B = 36'h000000000;
    parameter WRITE_MODE_A = "NO_CHANGE";
    parameter WRITE_MODE_B = "NO_CHANGE";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [31:0] CASDOUTA;
    output [31:0] CASDOUTB;
    output [3:0] CASDOUTPA;
    output [3:0] CASDOUTPB;
    output CASOUTDBITERR;
    output CASOUTSBITERR;
    output DBITERR;
    output [31:0] DOUTADOUT;
    output [31:0] DOUTBDOUT;
    output [3:0] DOUTPADOUTP;
    output [3:0] DOUTPBDOUTP;
    output [7:0] ECCPARITY;
    output [8:0] RDADDRECC;
    output SBITERR;
    input [14:0] ADDRARDADDR;
    input [14:0] ADDRBWRADDR;
    input ADDRENA;
    input ADDRENB;
    input CASDIMUXA;
    input CASDIMUXB;
    input [31:0] CASDINA;
    input [31:0] CASDINB;
    input [3:0] CASDINPA;
    input [3:0] CASDINPB;
    input CASDOMUXA;
    input CASDOMUXB;
    input CASDOMUXEN_A;
    input CASDOMUXEN_B;
    input CASINDBITERR;
    input CASINSBITERR;
    input CASOREGIMUXA;
    input CASOREGIMUXB;
    input CASOREGIMUXEN_A;
    input CASOREGIMUXEN_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKARDCLK_INVERTED" *)
    input CLKARDCLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKBWRCLK_INVERTED" *)
    input CLKBWRCLK;
    input [31:0] DINADIN;
    input [31:0] DINBDIN;
    input [3:0] DINPADINP;
    input [3:0] DINPBDINP;
    input ECCPIPECE;
    (* invertible_pin = "IS_ENARDEN_INVERTED" *)
    input ENARDEN;
    (* invertible_pin = "IS_ENBWREN_INVERTED" *)
    input ENBWREN;
    input INJECTDBITERR;
    input INJECTSBITERR;
    input REGCEAREGCE;
    input REGCEB;
    (* invertible_pin = "IS_RSTRAMARSTRAM_INVERTED" *)
    input RSTRAMARSTRAM;
    (* invertible_pin = "IS_RSTRAMB_INVERTED" *)
    input RSTRAMB;
    (* invertible_pin = "IS_RSTREGARSTREG_INVERTED" *)
    input RSTREGARSTREG;
    (* invertible_pin = "IS_RSTREGB_INVERTED" *)
    input RSTREGB;
    input SLEEP;
    input [3:0] WEA;
    input [7:0] WEBWE;
endmodule

module URAM288 (...);
    parameter integer AUTO_SLEEP_LATENCY = 8;
    parameter integer AVG_CONS_INACTIVE_CYCLES = 10;
    parameter BWE_MODE_A = "PARITY_INTERLEAVED";
    parameter BWE_MODE_B = "PARITY_INTERLEAVED";
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter EN_AUTO_SLEEP_MODE = "FALSE";
    parameter EN_ECC_RD_A = "FALSE";
    parameter EN_ECC_RD_B = "FALSE";
    parameter EN_ECC_WR_A = "FALSE";
    parameter EN_ECC_WR_B = "FALSE";
    parameter IREG_PRE_A = "FALSE";
    parameter IREG_PRE_B = "FALSE";
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_EN_A_INVERTED = 1'b0;
    parameter [0:0] IS_EN_B_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_A_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_B_INVERTED = 1'b0;
    parameter [0:0] IS_RST_A_INVERTED = 1'b0;
    parameter [0:0] IS_RST_B_INVERTED = 1'b0;
    parameter MATRIX_ID = "NONE";
    parameter integer NUM_UNIQUE_SELF_ADDR_A = 1;
    parameter integer NUM_UNIQUE_SELF_ADDR_B = 1;
    parameter integer NUM_URAM_IN_MATRIX = 1;
    parameter OREG_A = "FALSE";
    parameter OREG_B = "FALSE";
    parameter OREG_ECC_A = "FALSE";
    parameter OREG_ECC_B = "FALSE";
    parameter REG_CAS_A = "FALSE";
    parameter REG_CAS_B = "FALSE";
    parameter RST_MODE_A = "SYNC";
    parameter RST_MODE_B = "SYNC";
    parameter [10:0] SELF_ADDR_A = 11'h000;
    parameter [10:0] SELF_ADDR_B = 11'h000;
    parameter [10:0] SELF_MASK_A = 11'h7FF;
    parameter [10:0] SELF_MASK_B = 11'h7FF;
    parameter USE_EXT_CE_A = "FALSE";
    parameter USE_EXT_CE_B = "FALSE";
    output [22:0] CAS_OUT_ADDR_A;
    output [22:0] CAS_OUT_ADDR_B;
    output [8:0] CAS_OUT_BWE_A;
    output [8:0] CAS_OUT_BWE_B;
    output CAS_OUT_DBITERR_A;
    output CAS_OUT_DBITERR_B;
    output [71:0] CAS_OUT_DIN_A;
    output [71:0] CAS_OUT_DIN_B;
    output [71:0] CAS_OUT_DOUT_A;
    output [71:0] CAS_OUT_DOUT_B;
    output CAS_OUT_EN_A;
    output CAS_OUT_EN_B;
    output CAS_OUT_RDACCESS_A;
    output CAS_OUT_RDACCESS_B;
    output CAS_OUT_RDB_WR_A;
    output CAS_OUT_RDB_WR_B;
    output CAS_OUT_SBITERR_A;
    output CAS_OUT_SBITERR_B;
    output DBITERR_A;
    output DBITERR_B;
    output [71:0] DOUT_A;
    output [71:0] DOUT_B;
    output RDACCESS_A;
    output RDACCESS_B;
    output SBITERR_A;
    output SBITERR_B;
    input [22:0] ADDR_A;
    input [22:0] ADDR_B;
    input [8:0] BWE_A;
    input [8:0] BWE_B;
    input [22:0] CAS_IN_ADDR_A;
    input [22:0] CAS_IN_ADDR_B;
    input [8:0] CAS_IN_BWE_A;
    input [8:0] CAS_IN_BWE_B;
    input CAS_IN_DBITERR_A;
    input CAS_IN_DBITERR_B;
    input [71:0] CAS_IN_DIN_A;
    input [71:0] CAS_IN_DIN_B;
    input [71:0] CAS_IN_DOUT_A;
    input [71:0] CAS_IN_DOUT_B;
    input CAS_IN_EN_A;
    input CAS_IN_EN_B;
    input CAS_IN_RDACCESS_A;
    input CAS_IN_RDACCESS_B;
    input CAS_IN_RDB_WR_A;
    input CAS_IN_RDB_WR_B;
    input CAS_IN_SBITERR_A;
    input CAS_IN_SBITERR_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [71:0] DIN_A;
    input [71:0] DIN_B;
    (* invertible_pin = "IS_EN_A_INVERTED" *)
    input EN_A;
    (* invertible_pin = "IS_EN_B_INVERTED" *)
    input EN_B;
    input INJECT_DBITERR_A;
    input INJECT_DBITERR_B;
    input INJECT_SBITERR_A;
    input INJECT_SBITERR_B;
    input OREG_CE_A;
    input OREG_CE_B;
    input OREG_ECC_CE_A;
    input OREG_ECC_CE_B;
    (* invertible_pin = "IS_RDB_WR_A_INVERTED" *)
    input RDB_WR_A;
    (* invertible_pin = "IS_RDB_WR_B_INVERTED" *)
    input RDB_WR_B;
    (* invertible_pin = "IS_RST_A_INVERTED" *)
    input RST_A;
    (* invertible_pin = "IS_RST_B_INVERTED" *)
    input RST_B;
    input SLEEP;
endmodule

module URAM288_BASE (...);
    parameter integer AUTO_SLEEP_LATENCY = 8;
    parameter integer AVG_CONS_INACTIVE_CYCLES = 10;
    parameter BWE_MODE_A = "PARITY_INTERLEAVED";
    parameter BWE_MODE_B = "PARITY_INTERLEAVED";
    parameter EN_AUTO_SLEEP_MODE = "FALSE";
    parameter EN_ECC_RD_A = "FALSE";
    parameter EN_ECC_RD_B = "FALSE";
    parameter EN_ECC_WR_A = "FALSE";
    parameter EN_ECC_WR_B = "FALSE";
    parameter IREG_PRE_A = "FALSE";
    parameter IREG_PRE_B = "FALSE";
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_EN_A_INVERTED = 1'b0;
    parameter [0:0] IS_EN_B_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_A_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_B_INVERTED = 1'b0;
    parameter [0:0] IS_RST_A_INVERTED = 1'b0;
    parameter [0:0] IS_RST_B_INVERTED = 1'b0;
    parameter OREG_A = "FALSE";
    parameter OREG_B = "FALSE";
    parameter OREG_ECC_A = "FALSE";
    parameter OREG_ECC_B = "FALSE";
    parameter RST_MODE_A = "SYNC";
    parameter RST_MODE_B = "SYNC";
    parameter USE_EXT_CE_A = "FALSE";
    parameter USE_EXT_CE_B = "FALSE";
    output DBITERR_A;
    output DBITERR_B;
    output [71:0] DOUT_A;
    output [71:0] DOUT_B;
    output SBITERR_A;
    output SBITERR_B;
    input [22:0] ADDR_A;
    input [22:0] ADDR_B;
    input [8:0] BWE_A;
    input [8:0] BWE_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [71:0] DIN_A;
    input [71:0] DIN_B;
    (* invertible_pin = "IS_EN_A_INVERTED" *)
    input EN_A;
    (* invertible_pin = "IS_EN_B_INVERTED" *)
    input EN_B;
    input INJECT_DBITERR_A;
    input INJECT_DBITERR_B;
    input INJECT_SBITERR_A;
    input INJECT_SBITERR_B;
    input OREG_CE_A;
    input OREG_CE_B;
    input OREG_ECC_CE_A;
    input OREG_ECC_CE_B;
    (* invertible_pin = "IS_RDB_WR_A_INVERTED" *)
    input RDB_WR_A;
    (* invertible_pin = "IS_RDB_WR_B_INVERTED" *)
    input RDB_WR_B;
    (* invertible_pin = "IS_RST_A_INVERTED" *)
    input RST_A;
    (* invertible_pin = "IS_RST_B_INVERTED" *)
    input RST_B;
    input SLEEP;
endmodule

module DSP48E (...);
    parameter SIM_MODE = "SAFE";
    parameter integer ACASCREG = 1;
    parameter integer ALUMODEREG = 1;
    parameter integer AREG = 1;
    parameter AUTORESET_PATTERN_DETECT = "FALSE";
    parameter AUTORESET_PATTERN_DETECT_OPTINV = "MATCH";
    parameter A_INPUT = "DIRECT";
    parameter integer BCASCREG = 1;
    parameter integer BREG = 1;
    parameter B_INPUT = "DIRECT";
    parameter integer CARRYINREG = 1;
    parameter integer CARRYINSELREG = 1;
    parameter integer CREG = 1;
    parameter [47:0] MASK = 48'h3FFFFFFFFFFF;
    parameter integer MREG = 1;
    parameter integer MULTCARRYINREG = 1;
    parameter integer OPMODEREG = 1;
    parameter [47:0] PATTERN = 48'h000000000000;
    parameter integer PREG = 1;
    parameter SEL_MASK = "MASK";
    parameter SEL_PATTERN = "PATTERN";
    parameter SEL_ROUNDING_MASK = "SEL_MASK";
    parameter USE_MULT = "MULT_S";
    parameter USE_PATTERN_DETECT = "NO_PATDET";
    parameter USE_SIMD = "ONE48";
    output [29:0] ACOUT;
    output [17:0] BCOUT;
    output CARRYCASCOUT;
    output [3:0] CARRYOUT;
    output MULTSIGNOUT;
    output OVERFLOW;
    output [47:0] P;
    output PATTERNBDETECT;
    output PATTERNDETECT;
    output [47:0] PCOUT;
    output UNDERFLOW;
    input [29:0] A;
    input [29:0] ACIN;
    input [3:0] ALUMODE;
    input [17:0] B;
    input [17:0] BCIN;
    input [47:0] C;
    input CARRYCASCIN;
    input CARRYIN;
    input [2:0] CARRYINSEL;
    input CEA1;
    input CEA2;
    input CEALUMODE;
    input CEB1;
    input CEB2;
    input CEC;
    input CECARRYIN;
    input CECTRL;
    input CEM;
    input CEMULTCARRYIN;
    input CEP;
    (* clkbuf_sink *)
    input CLK;
    input MULTSIGNIN;
    input [6:0] OPMODE;
    input [47:0] PCIN;
    input RSTA;
    input RSTALLCARRYIN;
    input RSTALUMODE;
    input RSTB;
    input RSTC;
    input RSTCTRL;
    input RSTM;
    input RSTP;
endmodule

module DSP48E2 (...);
    parameter integer ACASCREG = 1;
    parameter integer ADREG = 1;
    parameter integer ALUMODEREG = 1;
    parameter AMULTSEL = "A";
    parameter integer AREG = 1;
    parameter AUTORESET_PATDET = "NO_RESET";
    parameter AUTORESET_PRIORITY = "RESET";
    parameter A_INPUT = "DIRECT";
    parameter integer BCASCREG = 1;
    parameter BMULTSEL = "B";
    parameter integer BREG = 1;
    parameter B_INPUT = "DIRECT";
    parameter integer CARRYINREG = 1;
    parameter integer CARRYINSELREG = 1;
    parameter integer CREG = 1;
    parameter integer DREG = 1;
    parameter integer INMODEREG = 1;
    parameter [3:0] IS_ALUMODE_INVERTED = 4'b0000;
    parameter [0:0] IS_CARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [4:0] IS_INMODE_INVERTED = 5'b00000;
    parameter [8:0] IS_OPMODE_INVERTED = 9'b000000000;
    parameter [0:0] IS_RSTALLCARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTALUMODE_INVERTED = 1'b0;
    parameter [0:0] IS_RSTA_INVERTED = 1'b0;
    parameter [0:0] IS_RSTB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTCTRL_INVERTED = 1'b0;
    parameter [0:0] IS_RSTC_INVERTED = 1'b0;
    parameter [0:0] IS_RSTD_INVERTED = 1'b0;
    parameter [0:0] IS_RSTINMODE_INVERTED = 1'b0;
    parameter [0:0] IS_RSTM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTP_INVERTED = 1'b0;
    parameter [47:0] MASK = 48'h3FFFFFFFFFFF;
    parameter integer MREG = 1;
    parameter integer OPMODEREG = 1;
    parameter [47:0] PATTERN = 48'h000000000000;
    parameter PREADDINSEL = "A";
    parameter integer PREG = 1;
    parameter [47:0] RND = 48'h000000000000;
    parameter SEL_MASK = "MASK";
    parameter SEL_PATTERN = "PATTERN";
    parameter USE_MULT = "MULTIPLY";
    parameter USE_PATTERN_DETECT = "NO_PATDET";
    parameter USE_SIMD = "ONE48";
    parameter USE_WIDEXOR = "FALSE";
    parameter XORSIMD = "XOR24_48_96";
    output [29:0] ACOUT;
    output [17:0] BCOUT;
    output CARRYCASCOUT;
    output [3:0] CARRYOUT;
    output MULTSIGNOUT;
    output OVERFLOW;
    output [47:0] P;
    output PATTERNBDETECT;
    output PATTERNDETECT;
    output [47:0] PCOUT;
    output UNDERFLOW;
    output [7:0] XOROUT;
    input [29:0] A;
    input [29:0] ACIN;
    (* invertible_pin = "IS_ALUMODE_INVERTED" *)
    input [3:0] ALUMODE;
    input [17:0] B;
    input [17:0] BCIN;
    input [47:0] C;
    input CARRYCASCIN;
    (* invertible_pin = "IS_CARRYIN_INVERTED" *)
    input CARRYIN;
    input [2:0] CARRYINSEL;
    input CEA1;
    input CEA2;
    input CEAD;
    input CEALUMODE;
    input CEB1;
    input CEB2;
    input CEC;
    input CECARRYIN;
    input CECTRL;
    input CED;
    input CEINMODE;
    input CEM;
    input CEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [26:0] D;
    (* invertible_pin = "IS_INMODE_INVERTED" *)
    input [4:0] INMODE;
    input MULTSIGNIN;
    (* invertible_pin = "IS_OPMODE_INVERTED" *)
    input [8:0] OPMODE;
    input [47:0] PCIN;
    (* invertible_pin = "IS_RSTA_INVERTED" *)
    input RSTA;
    (* invertible_pin = "IS_RSTALLCARRYIN_INVERTED" *)
    input RSTALLCARRYIN;
    (* invertible_pin = "IS_RSTALUMODE_INVERTED" *)
    input RSTALUMODE;
    (* invertible_pin = "IS_RSTB_INVERTED" *)
    input RSTB;
    (* invertible_pin = "IS_RSTC_INVERTED" *)
    input RSTC;
    (* invertible_pin = "IS_RSTCTRL_INVERTED" *)
    input RSTCTRL;
    (* invertible_pin = "IS_RSTD_INVERTED" *)
    input RSTD;
    (* invertible_pin = "IS_RSTINMODE_INVERTED" *)
    input RSTINMODE;
    (* invertible_pin = "IS_RSTM_INVERTED" *)
    input RSTM;
    (* invertible_pin = "IS_RSTP_INVERTED" *)
    input RSTP;
endmodule

module FDDRCPE (...);
    parameter INIT = 1'b0;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input D0;
    input D1;
    input CLR;
    input PRE;
    output Q;
endmodule

module FDDRRSE (...);
    parameter INIT = 1'b0;
    output Q;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input D0;
    input D1;
    input R;
    input S;
endmodule

module IFDDRCPE (...);
    output Q0;
    output Q1;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input CLR;
    (* iopad_external_pin *)
    input D;
    input PRE;
endmodule

module IFDDRRSE (...);
    output Q0;
    output Q1;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    (* iopad_external_pin *)
    input D;
    input R;
    input S;
endmodule

module OFDDRCPE (...);
    (* iopad_external_pin *)
    output Q;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input CLR;
    input D0;
    input D1;
    input PRE;
endmodule

module OFDDRRSE (...);
    (* iopad_external_pin *)
    output Q;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input D0;
    input D1;
    input R;
    input S;
endmodule

module OFDDRTCPE (...);
    (* iopad_external_pin *)
    output O;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input CLR;
    input D0;
    input D1;
    input PRE;
    input T;
endmodule

module OFDDRTRSE (...);
    (* iopad_external_pin *)
    output O;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input D0;
    input D1;
    input R;
    input S;
    input T;
endmodule

module IDDR2 (...);
    parameter DDR_ALIGNMENT = "NONE";
    parameter [0:0] INIT_Q0 = 1'b0;
    parameter [0:0] INIT_Q1 = 1'b0;
    parameter SRTYPE = "SYNC";
    output Q0;
    output Q1;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input D;
    input R;
    input S;
endmodule

module ODDR2 (...);
    parameter DDR_ALIGNMENT = "NONE";
    parameter [0:0] INIT = 1'b0;
    parameter SRTYPE = "SYNC";
    output Q;
    (* clkbuf_sink *)
    input C0;
    (* clkbuf_sink *)
    input C1;
    input CE;
    input D0;
    input D1;
    input R;
    input S;
endmodule

module IDDR (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter INIT_Q1 = 1'b0;
    parameter INIT_Q2 = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter SRTYPE = "SYNC";
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    input R;
    input S;
endmodule

module IDDR_2CLK (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter INIT_Q1 = 1'b0;
    parameter INIT_Q2 = 1'b0;
    parameter [0:0] IS_CB_INVERTED = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter SRTYPE = "SYNC";
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CB_INVERTED" *)
    input CB;
    input CE;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    input R;
    input S;
endmodule

module ODDR (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter INIT = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter SRTYPE = "SYNC";
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    (* invertible_pin = "IS_D1_INVERTED" *)
    input D1;
    (* invertible_pin = "IS_D2_INVERTED" *)
    input D2;
    input R;
    input S;
endmodule

(* keep *)
module IDELAYCTRL (...);
    parameter SIM_DEVICE = "7SERIES";
    output RDY;
    (* clkbuf_sink *)
    input REFCLK;
    input RST;
endmodule

module IDELAY (...);
    parameter IOBDELAY_TYPE = "DEFAULT";
    parameter integer IOBDELAY_VALUE = 0;
    output O;
    (* clkbuf_sink *)
    input C;
    input CE;
    input I;
    input INC;
    input RST;
endmodule

module ISERDES (...);
    parameter BITSLIP_ENABLE = "FALSE";
    parameter DATA_RATE = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter [0:0] INIT_Q1 = 1'b0;
    parameter [0:0] INIT_Q2 = 1'b0;
    parameter [0:0] INIT_Q3 = 1'b0;
    parameter [0:0] INIT_Q4 = 1'b0;
    parameter INTERFACE_TYPE = "MEMORY";
    parameter IOBDELAY = "NONE";
    parameter IOBDELAY_TYPE = "DEFAULT";
    parameter integer IOBDELAY_VALUE = 0;
    parameter integer NUM_CE = 2;
    parameter SERDES_MODE = "MASTER";
    parameter integer SIM_DELAY_D = 0;
    parameter integer SIM_SETUP_D_CLK = 0;
    parameter integer SIM_HOLD_D_CLK = 0;
    parameter [0:0] SRVAL_Q1 = 1'b0;
    parameter [0:0] SRVAL_Q2 = 1'b0;
    parameter [0:0] SRVAL_Q3 = 1'b0;
    parameter [0:0] SRVAL_Q4 = 1'b0;
    output O;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output SHIFTOUT1;
    output SHIFTOUT2;
    input BITSLIP;
    input CE1;
    input CE2;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    input D;
    input DLYCE;
    input DLYINC;
    input DLYRST;
    (* clkbuf_sink *)
    input OCLK;
    input REV;
    input SHIFTIN1;
    input SHIFTIN2;
    input SR;
endmodule

module OSERDES (...);
    parameter DATA_RATE_OQ = "DDR";
    parameter DATA_RATE_TQ = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter [0:0] INIT_OQ = 1'b0;
    parameter [0:0] INIT_TQ = 1'b0;
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_OQ = 1'b0;
    parameter [0:0] SRVAL_TQ = 1'b0;
    parameter integer TRISTATE_WIDTH = 4;
    output OQ;
    output SHIFTOUT1;
    output SHIFTOUT2;
    output TQ;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input OCE;
    input REV;
    input SHIFTIN1;
    input SHIFTIN2;
    input SR;
    input T1;
    input T2;
    input T3;
    input T4;
    input TCE;
endmodule

module IODELAY (...);
    parameter DELAY_SRC = "I";
    parameter HIGH_PERFORMANCE_MODE = "TRUE";
    parameter IDELAY_TYPE = "DEFAULT";
    parameter integer IDELAY_VALUE = 0;
    parameter integer ODELAY_VALUE = 0;
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    output DATAOUT;
    (* clkbuf_sink *)
    input C;
    input CE;
    input DATAIN;
    input IDATAIN;
    input INC;
    input ODATAIN;
    input RST;
    input T;
endmodule

module ISERDES_NODELAY (...);
    parameter BITSLIP_ENABLE = "FALSE";
    parameter DATA_RATE = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter INIT_Q1 = 1'b0;
    parameter INIT_Q2 = 1'b0;
    parameter INIT_Q3 = 1'b0;
    parameter INIT_Q4 = 1'b0;
    parameter INTERFACE_TYPE = "MEMORY";
    parameter integer NUM_CE = 2;
    parameter SERDES_MODE = "MASTER";
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output SHIFTOUT1;
    output SHIFTOUT2;
    input BITSLIP;
    input CE1;
    input CE2;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKB;
    (* clkbuf_sink *)
    input CLKDIV;
    input D;
    (* clkbuf_sink *)
    input OCLK;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
endmodule

module IODELAYE1 (...);
    parameter CINVCTRL_SEL = "FALSE";
    parameter DELAY_SRC = "I";
    parameter HIGH_PERFORMANCE_MODE = "FALSE";
    parameter IDELAY_TYPE = "DEFAULT";
    parameter integer IDELAY_VALUE = 0;
    parameter ODELAY_TYPE = "FIXED";
    parameter integer ODELAY_VALUE = 0;
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    output [4:0] CNTVALUEOUT;
    output DATAOUT;
    (* clkbuf_sink *)
    input C;
    input CE;
    input CINVCTRL;
    input CLKIN;
    input [4:0] CNTVALUEIN;
    input DATAIN;
    input IDATAIN;
    input INC;
    input ODATAIN;
    input RST;
    input T;
endmodule

module ISERDESE1 (...);
    parameter DATA_RATE = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter DYN_CLKDIV_INV_EN = "FALSE";
    parameter DYN_CLK_INV_EN = "FALSE";
    parameter [0:0] INIT_Q1 = 1'b0;
    parameter [0:0] INIT_Q2 = 1'b0;
    parameter [0:0] INIT_Q3 = 1'b0;
    parameter [0:0] INIT_Q4 = 1'b0;
    parameter INTERFACE_TYPE = "MEMORY";
    parameter integer NUM_CE = 2;
    parameter IOBDELAY = "NONE";
    parameter OFB_USED = "FALSE";
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_Q1 = 1'b0;
    parameter [0:0] SRVAL_Q2 = 1'b0;
    parameter [0:0] SRVAL_Q3 = 1'b0;
    parameter [0:0] SRVAL_Q4 = 1'b0;
    output O;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output SHIFTOUT1;
    output SHIFTOUT2;
    input BITSLIP;
    input CE1;
    input CE2;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKB;
    (* clkbuf_sink *)
    input CLKDIV;
    input D;
    input DDLY;
    input DYNCLKDIVSEL;
    input DYNCLKSEL;
    (* clkbuf_sink *)
    input OCLK;
    input OFB;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
endmodule

module OSERDESE1 (...);
    parameter DATA_RATE_OQ = "DDR";
    parameter DATA_RATE_TQ = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter integer DDR3_DATA = 1;
    parameter [0:0] INIT_OQ = 1'b0;
    parameter [0:0] INIT_TQ = 1'b0;
    parameter INTERFACE_TYPE = "DEFAULT";
    parameter integer ODELAY_USED = 0;
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_OQ = 1'b0;
    parameter [0:0] SRVAL_TQ = 1'b0;
    parameter integer TRISTATE_WIDTH = 4;
    output OCBEXTEND;
    output OFB;
    output OQ;
    output SHIFTOUT1;
    output SHIFTOUT2;
    output TFB;
    output TQ;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    input CLKPERF;
    input CLKPERFDELAY;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input OCE;
    input ODV;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
    input T1;
    input T2;
    input T3;
    input T4;
    input TCE;
    input WC;
endmodule

module IDELAYE2 (...);
    parameter CINVCTRL_SEL = "FALSE";
    parameter DELAY_SRC = "IDATAIN";
    parameter HIGH_PERFORMANCE_MODE = "FALSE";
    parameter IDELAY_TYPE = "FIXED";
    parameter integer IDELAY_VALUE = 0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_DATAIN_INVERTED = 1'b0;
    parameter [0:0] IS_IDATAIN_INVERTED = 1'b0;
    parameter PIPE_SEL = "FALSE";
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    parameter integer SIM_DELAY_D = 0;
    output [4:0] CNTVALUEOUT;
    output DATAOUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    input CINVCTRL;
    input [4:0] CNTVALUEIN;
    (* invertible_pin = "IS_DATAIN_INVERTED" *)
    input DATAIN;
    (* invertible_pin = "IS_IDATAIN_INVERTED" *)
    input IDATAIN;
    input INC;
    input LD;
    input LDPIPEEN;
    input REGRST;
endmodule

module ODELAYE2 (...);
    parameter CINVCTRL_SEL = "FALSE";
    parameter DELAY_SRC = "ODATAIN";
    parameter HIGH_PERFORMANCE_MODE = "FALSE";
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_ODATAIN_INVERTED = 1'b0;
    parameter ODELAY_TYPE = "FIXED";
    parameter integer ODELAY_VALUE = 0;
    parameter PIPE_SEL = "FALSE";
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    parameter integer SIM_DELAY_D = 0;
    output [4:0] CNTVALUEOUT;
    output DATAOUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    input CINVCTRL;
    input CLKIN;
    input [4:0] CNTVALUEIN;
    input INC;
    input LD;
    input LDPIPEEN;
    (* invertible_pin = "IS_ODATAIN_INVERTED" *)
    input ODATAIN;
    input REGRST;
endmodule

module ISERDESE2 (...);
    parameter DATA_RATE = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter DYN_CLKDIV_INV_EN = "FALSE";
    parameter DYN_CLK_INV_EN = "FALSE";
    parameter [0:0] INIT_Q1 = 1'b0;
    parameter [0:0] INIT_Q2 = 1'b0;
    parameter [0:0] INIT_Q3 = 1'b0;
    parameter [0:0] INIT_Q4 = 1'b0;
    parameter INTERFACE_TYPE = "MEMORY";
    parameter IOBDELAY = "NONE";
    parameter [0:0] IS_CLKB_INVERTED = 1'b0;
    parameter [0:0] IS_CLKDIVP_INVERTED = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter [0:0] IS_OCLKB_INVERTED = 1'b0;
    parameter [0:0] IS_OCLK_INVERTED = 1'b0;
    parameter integer NUM_CE = 2;
    parameter OFB_USED = "FALSE";
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_Q1 = 1'b0;
    parameter [0:0] SRVAL_Q2 = 1'b0;
    parameter [0:0] SRVAL_Q3 = 1'b0;
    parameter [0:0] SRVAL_Q4 = 1'b0;
    output O;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output Q7;
    output Q8;
    output SHIFTOUT1;
    output SHIFTOUT2;
    input BITSLIP;
    input CE1;
    input CE2;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKB_INVERTED" *)
    input CLKB;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIV_INVERTED" *)
    input CLKDIV;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIVP_INVERTED" *)
    input CLKDIVP;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    input DDLY;
    input DYNCLKDIVSEL;
    input DYNCLKSEL;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_OCLK_INVERTED" *)
    input OCLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_OCLKB_INVERTED" *)
    input OCLKB;
    input OFB;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
endmodule

module OSERDESE2 (...);
    parameter DATA_RATE_OQ = "DDR";
    parameter DATA_RATE_TQ = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter [0:0] INIT_OQ = 1'b0;
    parameter [0:0] INIT_TQ = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter [0:0] IS_D3_INVERTED = 1'b0;
    parameter [0:0] IS_D4_INVERTED = 1'b0;
    parameter [0:0] IS_D5_INVERTED = 1'b0;
    parameter [0:0] IS_D6_INVERTED = 1'b0;
    parameter [0:0] IS_D7_INVERTED = 1'b0;
    parameter [0:0] IS_D8_INVERTED = 1'b0;
    parameter [0:0] IS_T1_INVERTED = 1'b0;
    parameter [0:0] IS_T2_INVERTED = 1'b0;
    parameter [0:0] IS_T3_INVERTED = 1'b0;
    parameter [0:0] IS_T4_INVERTED = 1'b0;
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_OQ = 1'b0;
    parameter [0:0] SRVAL_TQ = 1'b0;
    parameter TBYTE_CTL = "FALSE";
    parameter TBYTE_SRC = "FALSE";
    parameter integer TRISTATE_WIDTH = 4;
    output OFB;
    output OQ;
    output SHIFTOUT1;
    output SHIFTOUT2;
    output TBYTEOUT;
    output TFB;
    output TQ;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIV_INVERTED" *)
    input CLKDIV;
    (* invertible_pin = "IS_D1_INVERTED" *)
    input D1;
    (* invertible_pin = "IS_D2_INVERTED" *)
    input D2;
    (* invertible_pin = "IS_D3_INVERTED" *)
    input D3;
    (* invertible_pin = "IS_D4_INVERTED" *)
    input D4;
    (* invertible_pin = "IS_D5_INVERTED" *)
    input D5;
    (* invertible_pin = "IS_D6_INVERTED" *)
    input D6;
    (* invertible_pin = "IS_D7_INVERTED" *)
    input D7;
    (* invertible_pin = "IS_D8_INVERTED" *)
    input D8;
    input OCE;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
    (* invertible_pin = "IS_T1_INVERTED" *)
    input T1;
    (* invertible_pin = "IS_T2_INVERTED" *)
    input T2;
    (* invertible_pin = "IS_T3_INVERTED" *)
    input T3;
    (* invertible_pin = "IS_T4_INVERTED" *)
    input T4;
    input TBYTEIN;
    input TCE;
endmodule

module PHASER_IN (...);
    parameter integer CLKOUT_DIV = 4;
    parameter DQS_BIAS_MODE = "FALSE";
    parameter EN_ISERDES_RST = "FALSE";
    parameter integer FINE_DELAY = 0;
    parameter FREQ_REF_DIV = "NONE";
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter integer SEL_CLK_OFFSET = 5;
    parameter SYNC_IN_DIV_RST = "FALSE";
    output FINEOVERFLOW;
    output ICLK;
    output ICLKDIV;
    output ISERDESRST;
    output RCLK;
    output [5:0] COUNTERREADVAL;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input DIVIDERST;
    input EDGEADV;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input SYNCIN;
    input SYSCLK;
    input [1:0] RANKSEL;
    input [5:0] COUNTERLOADVAL;
endmodule

module PHASER_IN_PHY (...);
    parameter BURST_MODE = "FALSE";
    parameter integer CLKOUT_DIV = 4;
    parameter [0:0] DQS_AUTO_RECAL = 1'b1;
    parameter DQS_BIAS_MODE = "FALSE";
    parameter [2:0] DQS_FIND_PATTERN = 3'b001;
    parameter integer FINE_DELAY = 0;
    parameter FREQ_REF_DIV = "NONE";
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter integer SEL_CLK_OFFSET = 5;
    parameter SYNC_IN_DIV_RST = "FALSE";
    parameter WR_CYCLES = "FALSE";
    output DQSFOUND;
    output DQSOUTOFRANGE;
    output FINEOVERFLOW;
    output ICLK;
    output ICLKDIV;
    output ISERDESRST;
    output PHASELOCKED;
    output RCLK;
    output WRENABLE;
    output [5:0] COUNTERREADVAL;
    input BURSTPENDINGPHY;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input RSTDQSFIND;
    input SYNCIN;
    input SYSCLK;
    input [1:0] ENCALIBPHY;
    input [1:0] RANKSELPHY;
    input [5:0] COUNTERLOADVAL;
endmodule

module PHASER_OUT (...);
    parameter integer CLKOUT_DIV = 4;
    parameter COARSE_BYPASS = "FALSE";
    parameter integer COARSE_DELAY = 0;
    parameter EN_OSERDES_RST = "FALSE";
    parameter integer FINE_DELAY = 0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OCLKDELAY_INV = "FALSE";
    parameter integer OCLK_DELAY = 0;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter [2:0] PO = 3'b000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter SYNC_IN_DIV_RST = "FALSE";
    output COARSEOVERFLOW;
    output FINEOVERFLOW;
    output OCLK;
    output OCLKDELAYED;
    output OCLKDIV;
    output OSERDESRST;
    output [8:0] COUNTERREADVAL;
    input COARSEENABLE;
    input COARSEINC;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input DIVIDERST;
    input EDGEADV;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input SELFINEOCLKDELAY;
    input SYNCIN;
    input SYSCLK;
    input [8:0] COUNTERLOADVAL;
endmodule

module PHASER_OUT_PHY (...);
    parameter integer CLKOUT_DIV = 4;
    parameter COARSE_BYPASS = "FALSE";
    parameter integer COARSE_DELAY = 0;
    parameter DATA_CTL_N = "FALSE";
    parameter DATA_RD_CYCLES = "FALSE";
    parameter integer FINE_DELAY = 0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OCLKDELAY_INV = "FALSE";
    parameter integer OCLK_DELAY = 0;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter [2:0] PO = 3'b000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter SYNC_IN_DIV_RST = "FALSE";
    output COARSEOVERFLOW;
    output FINEOVERFLOW;
    output OCLK;
    output OCLKDELAYED;
    output OCLKDIV;
    output OSERDESRST;
    output RDENABLE;
    output [1:0] CTSBUS;
    output [1:0] DQSBUS;
    output [1:0] DTSBUS;
    output [8:0] COUNTERREADVAL;
    input BURSTPENDINGPHY;
    input COARSEENABLE;
    input COARSEINC;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input SELFINEOCLKDELAY;
    input SYNCIN;
    input SYSCLK;
    input [1:0] ENCALIBPHY;
    input [8:0] COUNTERLOADVAL;
endmodule

module PHASER_REF (...);
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    output LOCKED;
    input CLKIN;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PHY_CONTROL (...);
    parameter integer AO_TOGGLE = 0;
    parameter [3:0] AO_WRLVL_EN = 4'b0000;
    parameter BURST_MODE = "FALSE";
    parameter integer CLK_RATIO = 1;
    parameter integer CMD_OFFSET = 0;
    parameter integer CO_DURATION = 0;
    parameter DATA_CTL_A_N = "FALSE";
    parameter DATA_CTL_B_N = "FALSE";
    parameter DATA_CTL_C_N = "FALSE";
    parameter DATA_CTL_D_N = "FALSE";
    parameter DISABLE_SEQ_MATCH = "TRUE";
    parameter integer DI_DURATION = 0;
    parameter integer DO_DURATION = 0;
    parameter integer EVENTS_DELAY = 63;
    parameter integer FOUR_WINDOW_CLOCKS = 63;
    parameter MULTI_REGION = "FALSE";
    parameter PHY_COUNT_ENABLE = "FALSE";
    parameter integer RD_CMD_OFFSET_0 = 0;
    parameter integer RD_CMD_OFFSET_1 = 00;
    parameter integer RD_CMD_OFFSET_2 = 0;
    parameter integer RD_CMD_OFFSET_3 = 0;
    parameter integer RD_DURATION_0 = 0;
    parameter integer RD_DURATION_1 = 0;
    parameter integer RD_DURATION_2 = 0;
    parameter integer RD_DURATION_3 = 0;
    parameter SYNC_MODE = "FALSE";
    parameter integer WR_CMD_OFFSET_0 = 0;
    parameter integer WR_CMD_OFFSET_1 = 0;
    parameter integer WR_CMD_OFFSET_2 = 0;
    parameter integer WR_CMD_OFFSET_3 = 0;
    parameter integer WR_DURATION_0 = 0;
    parameter integer WR_DURATION_1 = 0;
    parameter integer WR_DURATION_2 = 0;
    parameter integer WR_DURATION_3 = 0;
    output PHYCTLALMOSTFULL;
    output PHYCTLEMPTY;
    output PHYCTLFULL;
    output PHYCTLREADY;
    output [1:0] INRANKA;
    output [1:0] INRANKB;
    output [1:0] INRANKC;
    output [1:0] INRANKD;
    output [1:0] PCENABLECALIB;
    output [3:0] AUXOUTPUT;
    output [3:0] INBURSTPENDING;
    output [3:0] OUTBURSTPENDING;
    input MEMREFCLK;
    input PHYCLK;
    input PHYCTLMSTREMPTY;
    input PHYCTLWRENABLE;
    input PLLLOCK;
    input READCALIBENABLE;
    input REFDLLLOCK;
    input RESET;
    input SYNCIN;
    input WRITECALIBENABLE;
    input [31:0] PHYCTLWD;
endmodule

module IDDRE1 (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter [0:0] IS_CB_INVERTED = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CB_INVERTED" *)
    input CB;
    input D;
    input R;
endmodule

module ODDRE1 (...);
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter [0:0] SRVAL = 1'b0;
    output Q;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    (* invertible_pin = "IS_D1_INVERTED" *)
    input D1;
    (* invertible_pin = "IS_D2_INVERTED" *)
    input D2;
    input SR;
endmodule

module IDELAYE3 (...);
    parameter CASCADE = "NONE";
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_SRC = "IDATAIN";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter LOOPBACK = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output CASC_OUT;
    output [8:0] CNTVALUEOUT;
    output DATAOUT;
    input CASC_IN;
    input CASC_RETURN;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input DATAIN;
    input EN_VTC;
    input IDATAIN;
    input INC;
    input LOAD;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module ODELAYE3 (...);
    parameter CASCADE = "NONE";
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output CASC_OUT;
    output [8:0] CNTVALUEOUT;
    output DATAOUT;
    input CASC_IN;
    input CASC_RETURN;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input EN_VTC;
    input INC;
    input LOAD;
    input ODATAIN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module ISERDESE3 (...);
    parameter integer DATA_WIDTH = 8;
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter FIFO_ENABLE = "FALSE";
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter IDDR_MODE = "FALSE";
    parameter [0:0] IS_CLK_B_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output FIFO_EMPTY;
    output INTERNAL_DIVCLK;
    output [7:0] Q;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_B_INVERTED" *)
    input CLK_B;
    input D;
    (* clkbuf_sink *)
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module OSERDESE3 (...);
    parameter integer DATA_WIDTH = 8;
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter ODDR_MODE = "FALSE";
    parameter OSERDES_D_BYPASS = "FALSE";
    parameter OSERDES_T_BYPASS = "FALSE";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output OQ;
    output T_OUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIV_INVERTED" *)
    input CLKDIV;
    input [7:0] D;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input T;
endmodule

(* keep *)
module BITSLICE_CONTROL (...);
    parameter CTRL_CLK = "EXTERNAL";
    parameter DIV_MODE = "DIV2";
    parameter EN_CLK_TO_EXT_NORTH = "DISABLE";
    parameter EN_CLK_TO_EXT_SOUTH = "DISABLE";
    parameter EN_DYN_ODLY_MODE = "FALSE";
    parameter EN_OTHER_NCLK = "FALSE";
    parameter EN_OTHER_PCLK = "FALSE";
    parameter IDLY_VT_TRACK = "TRUE";
    parameter INV_RXCLK = "FALSE";
    parameter ODLY_VT_TRACK = "TRUE";
    parameter QDLY_VT_TRACK = "TRUE";
    parameter [5:0] READ_IDLE_COUNT = 6'h00;
    parameter REFCLK_SRC = "PLLCLK";
    parameter integer ROUNDING_FACTOR = 16;
    parameter RXGATE_EXTEND = "FALSE";
    parameter RX_CLK_PHASE_N = "SHIFT_0";
    parameter RX_CLK_PHASE_P = "SHIFT_0";
    parameter RX_GATING = "DISABLE";
    parameter SELF_CALIBRATE = "ENABLE";
    parameter SERIAL_MODE = "FALSE";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter SIM_SPEEDUP = "FAST";
    parameter real SIM_VERSION = 2.0;
    parameter TX_GATING = "DISABLE";
    output CLK_TO_EXT_NORTH;
    output CLK_TO_EXT_SOUTH;
    output DLY_RDY;
    output [6:0] DYN_DCI;
    output NCLK_NIBBLE_OUT;
    output PCLK_NIBBLE_OUT;
    output [15:0] RIU_RD_DATA;
    output RIU_VALID;
    output [39:0] RX_BIT_CTRL_OUT0;
    output [39:0] RX_BIT_CTRL_OUT1;
    output [39:0] RX_BIT_CTRL_OUT2;
    output [39:0] RX_BIT_CTRL_OUT3;
    output [39:0] RX_BIT_CTRL_OUT4;
    output [39:0] RX_BIT_CTRL_OUT5;
    output [39:0] RX_BIT_CTRL_OUT6;
    output [39:0] TX_BIT_CTRL_OUT0;
    output [39:0] TX_BIT_CTRL_OUT1;
    output [39:0] TX_BIT_CTRL_OUT2;
    output [39:0] TX_BIT_CTRL_OUT3;
    output [39:0] TX_BIT_CTRL_OUT4;
    output [39:0] TX_BIT_CTRL_OUT5;
    output [39:0] TX_BIT_CTRL_OUT6;
    output [39:0] TX_BIT_CTRL_OUT_TRI;
    output VTC_RDY;
    input CLK_FROM_EXT;
    input EN_VTC;
    input NCLK_NIBBLE_IN;
    input PCLK_NIBBLE_IN;
    input [3:0] PHY_RDCS0;
    input [3:0] PHY_RDCS1;
    input [3:0] PHY_RDEN;
    input [3:0] PHY_WRCS0;
    input [3:0] PHY_WRCS1;
    input PLL_CLK;
    input REFCLK;
    input [5:0] RIU_ADDR;
    input RIU_CLK;
    input RIU_NIBBLE_SEL;
    input [15:0] RIU_WR_DATA;
    input RIU_WR_EN;
    input RST;
    input [39:0] RX_BIT_CTRL_IN0;
    input [39:0] RX_BIT_CTRL_IN1;
    input [39:0] RX_BIT_CTRL_IN2;
    input [39:0] RX_BIT_CTRL_IN3;
    input [39:0] RX_BIT_CTRL_IN4;
    input [39:0] RX_BIT_CTRL_IN5;
    input [39:0] RX_BIT_CTRL_IN6;
    input [3:0] TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN0;
    input [39:0] TX_BIT_CTRL_IN1;
    input [39:0] TX_BIT_CTRL_IN2;
    input [39:0] TX_BIT_CTRL_IN3;
    input [39:0] TX_BIT_CTRL_IN4;
    input [39:0] TX_BIT_CTRL_IN5;
    input [39:0] TX_BIT_CTRL_IN6;
    input [39:0] TX_BIT_CTRL_IN_TRI;
endmodule

module RIU_OR (...);
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output [15:0] RIU_RD_DATA;
    output RIU_RD_VALID;
    input [15:0] RIU_RD_DATA_LOW;
    input [15:0] RIU_RD_DATA_UPP;
    input RIU_RD_VALID_LOW;
    input RIU_RD_VALID_UPP;
endmodule

module RX_BITSLICE (...);
    parameter CASCADE = "TRUE";
    parameter DATA_TYPE = "NONE";
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter integer DELAY_VALUE_EXT = 0;
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter [0:0] IS_CLK_EXT_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_EXT_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    parameter UPDATE_MODE_EXT = "ASYNC";
    output [8:0] CNTVALUEOUT;
    output [8:0] CNTVALUEOUT_EXT;
    output FIFO_EMPTY;
    output FIFO_WRCLK_OUT;
    output [7:0] Q;
    output [39:0] RX_BIT_CTRL_OUT;
    output [39:0] TX_BIT_CTRL_OUT;
    input CE;
    input CE_EXT;
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* invertible_pin = "IS_CLK_EXT_INVERTED" *)
    input CLK_EXT;
    input [8:0] CNTVALUEIN;
    input [8:0] CNTVALUEIN_EXT;
    input DATAIN;
    input EN_VTC;
    input EN_VTC_EXT;
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input INC;
    input INC_EXT;
    input LOAD;
    input LOAD_EXT;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RST_DLY_INVERTED" *)
    input RST_DLY;
    (* invertible_pin = "IS_RST_DLY_EXT_INVERTED" *)
    input RST_DLY_EXT;
    input [39:0] RX_BIT_CTRL_IN;
    input [39:0] TX_BIT_CTRL_IN;
endmodule

module RXTX_BITSLICE (...);
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_RX_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RX_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RX_RST_INVERTED = 1'b0;
    parameter [0:0] IS_TX_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_TX_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_TX_RST_INVERTED = 1'b0;
    parameter LOOPBACK = "FALSE";
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter ENABLE_PRE_EMPHASIS = "FALSE";
    parameter RX_DATA_TYPE = "NONE";
    parameter integer RX_DATA_WIDTH = 8;
    parameter RX_DELAY_FORMAT = "TIME";
    parameter RX_DELAY_TYPE = "FIXED";
    parameter integer RX_DELAY_VALUE = 0;
    parameter real RX_REFCLK_FREQUENCY = 300.0;
    parameter RX_UPDATE_MODE = "ASYNC";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter TBYTE_CTL = "TBYTE_IN";
    parameter integer TX_DATA_WIDTH = 8;
    parameter TX_DELAY_FORMAT = "TIME";
    parameter TX_DELAY_TYPE = "FIXED";
    parameter integer TX_DELAY_VALUE = 0;
    parameter TX_OUTPUT_PHASE_90 = "FALSE";
    parameter real TX_REFCLK_FREQUENCY = 300.0;
    parameter TX_UPDATE_MODE = "ASYNC";
    output FIFO_EMPTY;
    output FIFO_WRCLK_OUT;
    output O;
    output [7:0] Q;
    output [39:0] RX_BIT_CTRL_OUT;
    output [8:0] RX_CNTVALUEOUT;
    output [39:0] TX_BIT_CTRL_OUT;
    output [8:0] TX_CNTVALUEOUT;
    output T_OUT;
    input [7:0] D;
    input DATAIN;
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input [39:0] RX_BIT_CTRL_IN;
    input RX_CE;
    (* invertible_pin = "IS_RX_CLK_INVERTED" *)
    input RX_CLK;
    input [8:0] RX_CNTVALUEIN;
    input RX_EN_VTC;
    input RX_INC;
    input RX_LOAD;
    (* invertible_pin = "IS_RX_RST_INVERTED" *)
    input RX_RST;
    (* invertible_pin = "IS_RX_RST_DLY_INVERTED" *)
    input RX_RST_DLY;
    input T;
    input TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN;
    input TX_CE;
    (* invertible_pin = "IS_TX_CLK_INVERTED" *)
    input TX_CLK;
    input [8:0] TX_CNTVALUEIN;
    input TX_EN_VTC;
    input TX_INC;
    input TX_LOAD;
    (* invertible_pin = "IS_TX_RST_INVERTED" *)
    input TX_RST;
    (* invertible_pin = "IS_TX_RST_DLY_INVERTED" *)
    input TX_RST_DLY;
endmodule

module TX_BITSLICE (...);
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter ENABLE_PRE_EMPHASIS = "FALSE";
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter OUTPUT_PHASE_90 = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter TBYTE_CTL = "TBYTE_IN";
    parameter UPDATE_MODE = "ASYNC";
    output [8:0] CNTVALUEOUT;
    output O;
    output [39:0] RX_BIT_CTRL_OUT;
    output [39:0] TX_BIT_CTRL_OUT;
    output T_OUT;
    input CE;
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input [7:0] D;
    input EN_VTC;
    input INC;
    input LOAD;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RST_DLY_INVERTED" *)
    input RST_DLY;
    input [39:0] RX_BIT_CTRL_IN;
    input T;
    input TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN;
endmodule

module TX_BITSLICE_TRI (...);
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter OUTPUT_PHASE_90 = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output [39:0] BIT_CTRL_OUT;
    output [8:0] CNTVALUEOUT;
    output TRI_OUT;
    input [39:0] BIT_CTRL_IN;
    input CE;
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input EN_VTC;
    input INC;
    input LOAD;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RST_DLY_INVERTED" *)
    input RST_DLY;
endmodule

module IODELAY2 (...);
    parameter COUNTER_WRAPAROUND = "WRAPAROUND";
    parameter DATA_RATE = "SDR";
    parameter DELAY_SRC = "IO";
    parameter integer IDELAY2_VALUE = 0;
    parameter IDELAY_MODE = "NORMAL";
    parameter IDELAY_TYPE = "DEFAULT";
    parameter integer IDELAY_VALUE = 0;
    parameter integer ODELAY_VALUE = 0;
    parameter SERDES_MODE = "NONE";
    parameter integer SIM_TAPDELAY_VALUE = 75;
    output BUSY;
    output DATAOUT2;
    output DATAOUT;
    output DOUT;
    output TOUT;
    input CAL;
    input CE;
    (* clkbuf_sink *)
    input CLK;
    input IDATAIN;
    input INC;
    (* clkbuf_sink *)
    input IOCLK0;
    (* clkbuf_sink *)
    input IOCLK1;
    input ODATAIN;
    input RST;
    input T;
endmodule

module IODRP2 (...);
    parameter DATA_RATE = "SDR";
    parameter integer SIM_TAPDELAY_VALUE = 75;
    output DATAOUT2;
    output DATAOUT;
    output DOUT;
    output SDO;
    output TOUT;
    input ADD;
    input BKST;
    (* clkbuf_sink *)
    input CLK;
    input CS;
    input IDATAIN;
    (* clkbuf_sink *)
    input IOCLK0;
    (* clkbuf_sink *)
    input IOCLK1;
    input ODATAIN;
    input SDI;
    input T;
endmodule

module IODRP2_MCB (...);
    parameter DATA_RATE = "SDR";
    parameter integer IDELAY_VALUE = 0;
    parameter integer MCB_ADDRESS = 0;
    parameter integer ODELAY_VALUE = 0;
    parameter SERDES_MODE = "NONE";
    parameter integer SIM_TAPDELAY_VALUE = 75;
    output AUXSDO;
    output DATAOUT2;
    output DATAOUT;
    output DOUT;
    output DQSOUTN;
    output DQSOUTP;
    output SDO;
    output TOUT;
    input ADD;
    input AUXSDOIN;
    input BKST;
    (* clkbuf_sink *)
    input CLK;
    input CS;
    input IDATAIN;
    (* clkbuf_sink *)
    input IOCLK0;
    (* clkbuf_sink *)
    input IOCLK1;
    input MEMUPDATE;
    input ODATAIN;
    input SDI;
    input T;
    input [4:0] AUXADDR;
endmodule

module ISERDES2 (...);
    parameter BITSLIP_ENABLE = "FALSE";
    parameter DATA_RATE = "SDR";
    parameter integer DATA_WIDTH = 1;
    parameter INTERFACE_TYPE = "NETWORKING";
    parameter SERDES_MODE = "NONE";
    output CFB0;
    output CFB1;
    output DFB;
    output FABRICOUT;
    output INCDEC;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output SHIFTOUT;
    output VALID;
    input BITSLIP;
    input CE0;
    (* clkbuf_sink *)
    input CLK0;
    (* clkbuf_sink *)
    input CLK1;
    (* clkbuf_sink *)
    input CLKDIV;
    input D;
    input IOCE;
    input RST;
    input SHIFTIN;
endmodule

module OSERDES2 (...);
    parameter BYPASS_GCLK_FF = "FALSE";
    parameter DATA_RATE_OQ = "DDR";
    parameter DATA_RATE_OT = "DDR";
    parameter integer DATA_WIDTH = 2;
    parameter OUTPUT_MODE = "SINGLE_ENDED";
    parameter SERDES_MODE = "NONE";
    parameter integer TRAIN_PATTERN = 0;
    output OQ;
    output SHIFTOUT1;
    output SHIFTOUT2;
    output SHIFTOUT3;
    output SHIFTOUT4;
    output TQ;
    (* clkbuf_sink *)
    input CLK0;
    (* clkbuf_sink *)
    input CLK1;
    (* clkbuf_sink *)
    input CLKDIV;
    input D1;
    input D2;
    input D3;
    input D4;
    input IOCE;
    input OCE;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
    input SHIFTIN3;
    input SHIFTIN4;
    input T1;
    input T2;
    input T3;
    input T4;
    input TCE;
    input TRAIN;
endmodule

module IBUF_DLY_ADJ (...);
    parameter DELAY_OFFSET = "OFF";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    input [2:0] S;
endmodule

module IBUF_IBUFDISABLE (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
endmodule

module IBUF_INTERMDISABLE (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
endmodule

module IBUF_ANALOG (...);
    output O;
    (* iopad_external_pin *)
    input I;
endmodule

module IBUFE3 (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input OSC_EN;
    input VREF;
endmodule

module IBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IFD_DELAY_VALUE = "AUTO";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_DLY_ADJ (...);
    parameter DELAY_OFFSET = "OFF";
    parameter DIFF_TERM = "FALSE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input [2:0] S;
endmodule

module IBUFDS_IBUFDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
endmodule

module IBUFDS_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input INTERMDISABLE;
endmodule

module IBUFDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_DIFF_OUT_IBUFDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
endmodule

module IBUFDS_DIFF_OUT_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input INTERMDISABLE;
endmodule

module IBUFDSE3 (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input [3:0] OSC;
    input [1:0] OSC_EN;
endmodule

module IBUFDS_DPHY (...);
    parameter DIFF_TERM = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output HSRX_O;
    output LPRX_O_N;
    output LPRX_O_P;
    input HSRX_DISABLE;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input LPRX_DISABLE;
endmodule

module IBUFGDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter DIFF_TERM = "FALSE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFGDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IOBUF_DCIEN (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input T;
endmodule

module IOBUF_INTERMDISABLE (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
    input T;
endmodule

module IOBUFE3 (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    inout IO;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input OSC_EN;
    input T;
    input VREF;
endmodule

module IOBUFDS (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    output O;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input T;
endmodule

module IOBUFDS_DCIEN (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input T;
endmodule

module IOBUFDS_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter SLEW = "SLOW";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
    input T;
endmodule

module IOBUFDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input TM;
    input TS;
endmodule

module IOBUFDS_DIFF_OUT_DCIEN (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input TM;
    input TS;
endmodule

module IOBUFDS_DIFF_OUT_INTERMDISABLE (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SIM_DEVICE = "7SERIES";
    parameter USE_IBUFDISABLE = "TRUE";
    output O;
    output OB;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input I;
    input IBUFDISABLE;
    input INTERMDISABLE;
    input TM;
    input TS;
endmodule

module IOBUFDSE3 (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    parameter USE_IBUFDISABLE = "FALSE";
    output O;
    (* iopad_external_pin *)
    inout IO;
    (* iopad_external_pin *)
    inout IOB;
    input DCITERMDISABLE;
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input [1:0] OSC_EN;
    input T;
endmodule

module OBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
endmodule

module OBUFDS_DPHY (...);
    parameter IOSTANDARD = "DEFAULT";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input HSTX_I;
    input HSTX_T;
    input LPTX_I_N;
    input LPTX_I_P;
    input LPTX_T;
endmodule

module OBUFTDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
    input T;
endmodule

module KEEPER (...);
    inout O;
endmodule

module PULLDOWN (...);
    output O;
endmodule

module PULLUP (...);
    output O;
endmodule

(* keep *)
module DCIRESET (...);
    output LOCKED;
    input RST;
endmodule

module HPIO_VREF (...);
    parameter VREF_CNTR = "OFF";
    output VREF;
    input [6:0] FABRIC_VREF_TUNE;
endmodule

module BUFGCE (...);
    parameter CE_TYPE = "SYNC";
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter STARTUP_SYNC = "FALSE";
    (* clkbuf_driver *)
    output O;
    (* invertible_pin = "IS_CE_INVERTED" *)
    input CE;
    (* invertible_pin = "IS_I_INVERTED" *)
    input I;
endmodule

module BUFGCE_1 (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input I;
endmodule

module BUFGMUX (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_1 (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_CTRL (...);
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_VIRTEX4 (...);
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFG_GT (...);
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter STARTUP_SYNC = "FALSE";
    (* clkbuf_driver *)
    output O;
    input CE;
    input CEMASK;
    input CLR;
    input CLRMASK;
    input [2:0] DIV;
    input I;
endmodule

module BUFG_GT_SYNC (...);
    output CESYNC;
    output CLRSYNC;
    input CE;
    input CLK;
    input CLR;
endmodule

module BUFG_PS (...);
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter STARTUP_SYNC = "FALSE";
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFGCE_DIV (...);
    parameter integer BUFGCE_DIVIDE = 1;
    parameter CE_TYPE = "SYNC";
    parameter HARDSYNC_CLR = "FALSE";
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter STARTUP_SYNC = "FALSE";
    (* clkbuf_driver *)
    output O;
    (* invertible_pin = "IS_CE_INVERTED" *)
    input CE;
    (* invertible_pin = "IS_CLR_INVERTED" *)
    input CLR;
    (* invertible_pin = "IS_I_INVERTED" *)
    input I;
endmodule

module BUFH (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFIO2 (...);
    parameter DIVIDE_BYPASS = "TRUE";
    parameter integer DIVIDE = 1;
    parameter I_INVERT = "FALSE";
    parameter USE_DOUBLER = "FALSE";
    (* clkbuf_driver *)
    output DIVCLK;
    (* clkbuf_driver *)
    output IOCLK;
    output SERDESSTROBE;
    input I;
endmodule

module BUFIO2_2CLK (...);
    parameter integer DIVIDE = 2;
    (* clkbuf_driver *)
    output DIVCLK;
    (* clkbuf_driver *)
    output IOCLK;
    output SERDESSTROBE;
    input I;
    input IB;
endmodule

module BUFIO2FB (...);
    parameter DIVIDE_BYPASS = "TRUE";
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFPLL (...);
    parameter integer DIVIDE = 1;
    parameter ENABLE_SYNC = "TRUE";
    (* clkbuf_driver *)
    output IOCLK;
    output LOCK;
    output SERDESSTROBE;
    input GCLK;
    input LOCKED;
    input PLLIN;
endmodule

module BUFPLL_MCB (...);
    parameter integer DIVIDE = 2;
    parameter LOCK_SRC = "LOCK_TO_0";
    (* clkbuf_driver *)
    output IOCLK0;
    (* clkbuf_driver *)
    output IOCLK1;
    output LOCK;
    output SERDESSTROBE0;
    output SERDESSTROBE1;
    input GCLK;
    input LOCKED;
    input PLLIN0;
    input PLLIN1;
endmodule

module BUFIO (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFIODQS (...);
    parameter DQSMASK_ENABLE = "FALSE";
    (* clkbuf_driver *)
    output O;
    input DQSMASK;
    input I;
endmodule

module BUFR (...);
    parameter BUFR_DIVIDE = "BYPASS";
    parameter SIM_DEVICE = "7SERIES";
    (* clkbuf_driver *)
    output O;
    input CE;
    input CLR;
    input I;
endmodule

module BUFMR (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFMRCE (...);
    parameter CE_TYPE = "SYNC";
    parameter integer INIT_OUT = 0;
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    (* invertible_pin = "IS_CE_INVERTED" *)
    input CE;
    input I;
endmodule

module DCM (...);
    parameter real CLKDV_DIVIDE = 2.0;
    parameter integer CLKFX_DIVIDE = 1;
    parameter integer CLKFX_MULTIPLY = 4;
    parameter CLKIN_DIVIDE_BY_2 = "FALSE";
    parameter real CLKIN_PERIOD = 10.0;
    parameter CLKOUT_PHASE_SHIFT = "NONE";
    parameter CLK_FEEDBACK = "1X";
    parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
    parameter DFS_FREQUENCY_MODE = "LOW";
    parameter DLL_FREQUENCY_MODE = "LOW";
    parameter DSS_MODE = "NONE";
    parameter DUTY_CYCLE_CORRECTION = "TRUE";
    parameter [15:0] FACTORY_JF = 16'hC080;
    parameter integer PHASE_SHIFT = 0;
    parameter SIM_MODE = "SAFE";
    parameter STARTUP_WAIT = "FALSE";
    input CLKFB;
    input CLKIN;
    input DSSEN;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input RST;
    output CLK0;
    output CLK180;
    output CLK270;
    output CLK2X;
    output CLK2X180;
    output CLK90;
    output CLKDV;
    output CLKFX;
    output CLKFX180;
    output LOCKED;
    output PSDONE;
    output [7:0] STATUS;
endmodule

module DCM_SP (...);
    parameter real CLKDV_DIVIDE = 2.0;
    parameter integer CLKFX_DIVIDE = 1;
    parameter integer CLKFX_MULTIPLY = 4;
    parameter CLKIN_DIVIDE_BY_2 = "FALSE";
    parameter real CLKIN_PERIOD = 10.0;
    parameter CLKOUT_PHASE_SHIFT = "NONE";
    parameter CLK_FEEDBACK = "1X";
    parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
    parameter DFS_FREQUENCY_MODE = "LOW";
    parameter DLL_FREQUENCY_MODE = "LOW";
    parameter DSS_MODE = "NONE";
    parameter DUTY_CYCLE_CORRECTION = "TRUE";
    parameter FACTORY_JF = 16'hC080;
    parameter integer PHASE_SHIFT = 0;
    parameter STARTUP_WAIT = "FALSE";
    input CLKFB;
    input CLKIN;
    input DSSEN;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input RST;
    output CLK0;
    output CLK180;
    output CLK270;
    output CLK2X;
    output CLK2X180;
    output CLK90;
    output CLKDV;
    output CLKFX;
    output CLKFX180;
    output LOCKED;
    output PSDONE;
    output [7:0] STATUS;
endmodule

module DCM_CLKGEN (...);
    parameter SPREAD_SPECTRUM = "NONE";
    parameter STARTUP_WAIT = "FALSE";
    parameter integer CLKFXDV_DIVIDE = 2;
    parameter integer CLKFX_DIVIDE = 1;
    parameter integer CLKFX_MULTIPLY = 4;
    parameter real CLKFX_MD_MAX = 0.0;
    parameter real CLKIN_PERIOD = 0.0;
    output CLKFX180;
    output CLKFX;
    output CLKFXDV;
    output LOCKED;
    output PROGDONE;
    output [2:1] STATUS;
    input CLKIN;
    input FREEZEDCM;
    input PROGCLK;
    input PROGDATA;
    input PROGEN;
    input RST;
endmodule

module DCM_ADV (...);
    parameter real CLKDV_DIVIDE = 2.0;
    parameter integer CLKFX_DIVIDE = 1;
    parameter integer CLKFX_MULTIPLY = 4;
    parameter CLKIN_DIVIDE_BY_2 = "FALSE";
    parameter real CLKIN_PERIOD = 10.0;
    parameter CLKOUT_PHASE_SHIFT = "NONE";
    parameter CLK_FEEDBACK = "1X";
    parameter DCM_AUTOCALIBRATION = "TRUE";
    parameter DCM_PERFORMANCE_MODE = "MAX_SPEED";
    parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
    parameter DFS_FREQUENCY_MODE = "LOW";
    parameter DLL_FREQUENCY_MODE = "LOW";
    parameter DUTY_CYCLE_CORRECTION = "TRUE";
    parameter FACTORY_JF = 16'hF0F0;
    parameter integer PHASE_SHIFT = 0;
    parameter SIM_DEVICE ="VIRTEX4";
    parameter STARTUP_WAIT = "FALSE";
    output CLK0;
    output CLK180;
    output CLK270;
    output CLK2X180;
    output CLK2X;
    output CLK90;
    output CLKDV;
    output CLKFX180;
    output CLKFX;
    output DRDY;
    output LOCKED;
    output PSDONE;
    output [15:0] DO;
    input CLKFB;
    input CLKIN;
    input DCLK;
    input DEN;
    input DWE;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input RST;
    input [15:0] DI;
    input [6:0] DADDR;
endmodule

module DCM_BASE (...);
    parameter real CLKDV_DIVIDE = 2.0;
    parameter integer CLKFX_DIVIDE = 1;
    parameter integer CLKFX_MULTIPLY = 4;
    parameter CLKIN_DIVIDE_BY_2 = "FALSE";
    parameter real CLKIN_PERIOD = 10.0;
    parameter CLKOUT_PHASE_SHIFT = "NONE";
    parameter CLK_FEEDBACK = "1X";
    parameter DCM_AUTOCALIBRATION = "TRUE";
    parameter DCM_PERFORMANCE_MODE = "MAX_SPEED";
    parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
    parameter DFS_FREQUENCY_MODE = "LOW";
    parameter DLL_FREQUENCY_MODE = "LOW";
    parameter DUTY_CYCLE_CORRECTION = "TRUE";
    parameter [15:0] FACTORY_JF = 16'hF0F0;
    parameter integer PHASE_SHIFT = 0;
    parameter STARTUP_WAIT = "FALSE";
    output CLK0;
    output CLK180;
    output CLK270;
    output CLK2X180;
    output CLK2X;
    output CLK90;
    output CLKDV;
    output CLKFX180;
    output CLKFX;
    output LOCKED;
    input CLKFB;
    input CLKIN;
    input RST;
endmodule

module DCM_PS (...);
    parameter real CLKDV_DIVIDE = 2.0;
    parameter integer CLKFX_DIVIDE = 1;
    parameter integer CLKFX_MULTIPLY = 4;
    parameter CLKIN_DIVIDE_BY_2 = "FALSE";
    parameter real CLKIN_PERIOD = 10.0;
    parameter CLKOUT_PHASE_SHIFT = "NONE";
    parameter CLK_FEEDBACK = "1X";
    parameter DCM_AUTOCALIBRATION = "TRUE";
    parameter DCM_PERFORMANCE_MODE = "MAX_SPEED";
    parameter DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS";
    parameter DFS_FREQUENCY_MODE = "LOW";
    parameter DLL_FREQUENCY_MODE = "LOW";
    parameter DUTY_CYCLE_CORRECTION = "TRUE";
    parameter [15:0] FACTORY_JF = 16'hF0F0;
    parameter integer PHASE_SHIFT = 0;
    parameter STARTUP_WAIT = "FALSE";
    output CLK0;
    output CLK180;
    output CLK270;
    output CLK2X180;
    output CLK2X;
    output CLK90;
    output CLKDV;
    output CLKFX180;
    output CLKFX;
    output LOCKED;
    output PSDONE;
    output [15:0] DO;
    input CLKFB;
    input CLKIN;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input RST;
endmodule

module PMCD (...);
    parameter EN_REL = "FALSE";
    parameter RST_DEASSERT_CLK = "CLKA";
    output CLKA1;
    output CLKA1D2;
    output CLKA1D4;
    output CLKA1D8;
    output CLKB1;
    output CLKC1;
    output CLKD1;
    input CLKA;
    input CLKB;
    input CLKC;
    input CLKD;
    input REL;
    input RST;
endmodule

module PLL_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter CLK_FEEDBACK = "CLKFBOUT";
    parameter CLKFBOUT_DESKEW_ADJUST = "NONE";
    parameter CLKOUT0_DESKEW_ADJUST = "NONE";
    parameter CLKOUT1_DESKEW_ADJUST = "NONE";
    parameter CLKOUT2_DESKEW_ADJUST = "NONE";
    parameter CLKOUT3_DESKEW_ADJUST = "NONE";
    parameter CLKOUT4_DESKEW_ADJUST = "NONE";
    parameter CLKOUT5_DESKEW_ADJUST = "NONE";
    parameter integer CLKFBOUT_MULT = 1;
    parameter real CLKFBOUT_PHASE = 0.0;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.5;
    parameter real CLKOUT0_PHASE = 0.0;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.5;
    parameter real CLKOUT1_PHASE = 0.0;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.5;
    parameter real CLKOUT2_PHASE = 0.0;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.5;
    parameter real CLKOUT3_PHASE = 0.0;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.5;
    parameter real CLKOUT4_PHASE = 0.0;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.5;
    parameter real CLKOUT5_PHASE = 0.0;
    parameter COMPENSATION = "SYSTEM_SYNCHRONOUS";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter EN_REL = "FALSE";
    parameter PLL_PMCD_MODE = "FALSE";
    parameter real REF_JITTER = 0.100;
    parameter RESET_ON_LOSS_OF_LOCK = "FALSE";
    parameter RST_DEASSERT_CLK = "CLKIN1";
    parameter SIM_DEVICE = "VIRTEX5";
    parameter real VCOCLK_FREQ_MAX = 1440.0;
    parameter real VCOCLK_FREQ_MIN = 400.0;
    parameter real CLKIN_FREQ_MAX = 710.0;
    parameter real CLKIN_FREQ_MIN = 19.0;
    parameter real CLKPFD_FREQ_MAX = 550.0;
    parameter real CLKPFD_FREQ_MIN = 19.0;
    output CLKFBDCM;
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT1;
    output CLKOUT2;
    output CLKOUT3;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUTDCM0;
    output CLKOUTDCM1;
    output CLKOUTDCM2;
    output CLKOUTDCM3;
    output CLKOUTDCM4;
    output CLKOUTDCM5;
    output DRDY;
    output LOCKED;
    output [15:0] DO;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    input CLKINSEL;
    input DCLK;
    input DEN;
    input DWE;
    input REL;
    input RST;
    input [15:0] DI;
    input [4:0] DADDR;
endmodule

module PLL_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter integer CLKFBOUT_MULT = 1;
    parameter real CLKFBOUT_PHASE = 0.0;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.5;
    parameter real CLKOUT0_PHASE = 0.0;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.5;
    parameter real CLKOUT1_PHASE = 0.0;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.5;
    parameter real CLKOUT2_PHASE = 0.0;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.5;
    parameter real CLKOUT3_PHASE = 0.0;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.5;
    parameter real CLKOUT4_PHASE = 0.0;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.5;
    parameter real CLKOUT5_PHASE = 0.0;
    parameter CLK_FEEDBACK = "CLKFBOUT";
    parameter COMPENSATION = "SYSTEM_SYNCHRONOUS";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER = 0.100;
    parameter RESET_ON_LOSS_OF_LOCK = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT1;
    output CLKOUT2;
    output CLKOUT3;
    output CLKOUT4;
    output CLKOUT5;
    output LOCKED;
    input CLKFBIN;
    input CLKIN;
    input RST;
endmodule

module MMCM_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter CLOCK_HOLD = "FALSE";
    parameter COMPENSATION = "ZHOLD";
    parameter STARTUP_WAIT = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter real VCOCLK_FREQ_MAX = 1600.0;
    parameter real VCOCLK_FREQ_MIN = 600.0;
    parameter real CLKIN_FREQ_MAX = 800.0;
    parameter real CLKIN_FREQ_MIN = 10.0;
    parameter real CLKPFD_FREQ_MAX = 550.0;
    parameter real CLKPFD_FREQ_MIN = 10.0;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output DRDY;
    output LOCKED;
    output PSDONE;
    output [15:0] DO;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    input CLKINSEL;
    input DCLK;
    input DEN;
    input DWE;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input PWRDWN;
    input RST;
    input [15:0] DI;
    input [6:0] DADDR;
endmodule

module MMCM_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLOCK_HOLD = "FALSE";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module MMCME2_ADV (...);
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter COMPENSATION = "ZHOLD";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    (* invertible_pin = "IS_PSEN_INVERTED" *)
    input PSEN;
    (* invertible_pin = "IS_PSINCDEC_INVERTED" *)
    input PSINCDEC;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME2_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module PLLE2_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter COMPENSATION = "ZHOLD";
    parameter STARTUP_WAIT = "FALSE";
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter real VCOCLK_FREQ_MAX = 2133.000;
    parameter real VCOCLK_FREQ_MIN = 800.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 19.000;
    parameter real CLKPFD_FREQ_MAX = 550.0;
    parameter real CLKPFD_FREQ_MIN = 19.0;
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT1;
    output CLKOUT2;
    output CLKOUT3;
    output CLKOUT4;
    output CLKOUT5;
    output DRDY;
    output LOCKED;
    output [15:0] DO;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input DCLK;
    input DEN;
    input DWE;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input [15:0] DI;
    input [6:0] DADDR;
endmodule

module PLLE2_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT1;
    output CLKOUT2;
    output CLKOUT3;
    output CLKOUT4;
    output CLKOUT5;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module MMCME3_ADV (...);
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN2_INVERTED = 1'b0;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    output CDDCDONE;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CDDCREQ;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_CLKIN2_INVERTED" *)
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    (* invertible_pin = "IS_PSEN_INVERTED" *)
    input PSEN;
    (* invertible_pin = "IS_PSINCDEC_INVERTED" *)
    input PSINCDEC;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME3_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE3_ADV (...);
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 70.000;
    parameter real CLKPFD_FREQ_MAX = 667.500;
    parameter real CLKPFD_FREQ_MIN = 70.000;
    parameter real VCOCLK_FREQ_MAX = 1335.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE3_BASE (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME4_ADV (...);
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 800.000;
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN2_INVERTED = 1'b0;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    output CDDCDONE;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CDDCREQ;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_CLKIN2_INVERTED" *)
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    (* invertible_pin = "IS_PSEN_INVERTED" *)
    input PSEN;
    (* invertible_pin = "IS_PSINCDEC_INVERTED" *)
    input PSINCDEC;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME4_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE4_ADV (...);
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 70.000;
    parameter real CLKPFD_FREQ_MAX = 667.500;
    parameter real CLKPFD_FREQ_MIN = 70.000;
    parameter real VCOCLK_FREQ_MAX = 1500.000;
    parameter real VCOCLK_FREQ_MIN = 750.000;
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE4_BASE (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module BUFT (...);
    output O;
    input I;
    input T;
endmodule

module IN_FIFO (...);
    parameter integer ALMOST_EMPTY_VALUE = 1;
    parameter integer ALMOST_FULL_VALUE = 1;
    parameter ARRAY_MODE = "ARRAY_MODE_4_X_8";
    parameter SYNCHRONOUS_MODE = "FALSE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output EMPTY;
    output FULL;
    output [7:0] Q0;
    output [7:0] Q1;
    output [7:0] Q2;
    output [7:0] Q3;
    output [7:0] Q4;
    output [7:0] Q5;
    output [7:0] Q6;
    output [7:0] Q7;
    output [7:0] Q8;
    output [7:0] Q9;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RESET;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [3:0] D0;
    input [3:0] D1;
    input [3:0] D2;
    input [3:0] D3;
    input [3:0] D4;
    input [3:0] D7;
    input [3:0] D8;
    input [3:0] D9;
    input [7:0] D5;
    input [7:0] D6;
endmodule

module OUT_FIFO (...);
    parameter integer ALMOST_EMPTY_VALUE = 1;
    parameter integer ALMOST_FULL_VALUE = 1;
    parameter ARRAY_MODE = "ARRAY_MODE_8_X_4";
    parameter OUTPUT_DISABLE = "FALSE";
    parameter SYNCHRONOUS_MODE = "FALSE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output EMPTY;
    output FULL;
    output [3:0] Q0;
    output [3:0] Q1;
    output [3:0] Q2;
    output [3:0] Q3;
    output [3:0] Q4;
    output [3:0] Q7;
    output [3:0] Q8;
    output [3:0] Q9;
    output [7:0] Q5;
    output [7:0] Q6;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RESET;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [7:0] D0;
    input [7:0] D1;
    input [7:0] D2;
    input [7:0] D3;
    input [7:0] D4;
    input [7:0] D5;
    input [7:0] D6;
    input [7:0] D7;
    input [7:0] D8;
    input [7:0] D9;
endmodule

module HARD_SYNC (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter integer LATENCY = 2;
    output DOUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input DIN;
endmodule

(* keep *)
module STARTUP_SPARTAN3 (...);
    input CLK;
    input GSR;
    input GTS;
endmodule

(* keep *)
module STARTUP_SPARTAN3E (...);
    input CLK;
    input GSR;
    input GTS;
    input MBT;
endmodule

(* keep *)
module STARTUP_SPARTAN3A (...);
    input CLK;
    input GSR;
    input GTS;
endmodule

(* keep *)
module STARTUP_SPARTAN6 (...);
    output CFGCLK;
    output CFGMCLK;
    output EOS;
    input CLK;
    input GSR;
    input GTS;
    input KEYCLEARB;
endmodule

(* keep *)
module STARTUP_VIRTEX4 (...);
    output EOS;
    input CLK;
    input GSR;
    input GTS;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUP_VIRTEX5 (...);
    output CFGCLK;
    output CFGMCLK;
    output DINSPI;
    output EOS;
    output TCKSPI;
    input CLK;
    input GSR;
    input GTS;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUP_VIRTEX6 (...);
    parameter PROG_USR = "FALSE";
    output CFGCLK;
    output CFGMCLK;
    output DINSPI;
    output EOS;
    output PREQ;
    output TCKSPI;
    input CLK;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUPE2 (...);
    parameter PROG_USR = "FALSE";
    parameter real SIM_CCLK_FREQ = 0.0;
    output CFGCLK;
    output CFGMCLK;
    output EOS;
    output PREQ;
    input CLK;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUPE3 (...);
    parameter PROG_USR = "FALSE";
    parameter real SIM_CCLK_FREQ = 0.0;
    output CFGCLK;
    output CFGMCLK;
    output [3:0] DI;
    output EOS;
    output PREQ;
    input [3:0] DO;
    input [3:0] DTS;
    input FCSBO;
    input FCSBTS;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module CAPTURE_SPARTAN3 (...);
    parameter ONESHOT = "FALSE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTURE_SPARTAN3A (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTURE_VIRTEX4 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTURE_VIRTEX5 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTURE_VIRTEX6 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTUREE2 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module ICAP_SPARTAN3A (...);
    output BUSY;
    output [7:0] O;
    input CE;
    input CLK;
    input WRITE;
    input [7:0] I;
endmodule

(* keep *)
module ICAP_SPARTAN6 (...);
    parameter DEVICE_ID = 32'h04000093;
    parameter SIM_CFG_FILE_NAME = "NONE";
    output BUSY;
    output [15:0] O;
    input CLK;
    input CE;
    input WRITE;
    input [15:0] I;
endmodule

(* keep *)
module ICAP_VIRTEX4 (...);
    parameter ICAP_WIDTH = "X8";
    output BUSY;
    output [31:0] O;
    input CE;
    input CLK;
    input WRITE;
    input [31:0] I;
endmodule

(* keep *)
module ICAP_VIRTEX5 (...);
    parameter ICAP_WIDTH = "X8";
    output BUSY;
    output [31:0] O;
    input CE;
    input CLK;
    input WRITE;
    input [31:0] I;
endmodule

(* keep *)
module ICAP_VIRTEX6 (...);
    parameter [31:0] DEVICE_ID = 32'h04244093;
    parameter ICAP_WIDTH = "X8";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output BUSY;
    output [31:0] O;
    input CLK;
    input CSB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module ICAPE2 (...);
    parameter [31:0] DEVICE_ID = 32'h04244093;
    parameter ICAP_WIDTH = "X32";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output [31:0] O;
    input CLK;
    input CSIB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module ICAPE3 (...);
    parameter [31:0] DEVICE_ID = 32'h03628093;
    parameter ICAP_AUTO_SWITCH = "DISABLE";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output AVAIL;
    output [31:0] O;
    output PRDONE;
    output PRERROR;
    input CLK;
    input CSIB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module BSCAN_SPARTAN3 (...);
    output CAPTURE;
    output DRCK1;
    output DRCK2;
    output RESET;
    output SEL1;
    output SEL2;
    output SHIFT;
    output TDI;
    output UPDATE;
    input TDO1;
    input TDO2;
endmodule

(* keep *)
module BSCAN_SPARTAN3A (...);
    output CAPTURE;
    output DRCK1;
    output DRCK2;
    output RESET;
    output SEL1;
    output SEL2;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO1;
    input TDO2;
endmodule

(* keep *)
module BSCAN_SPARTAN6 (...);
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCAN_VIRTEX4 (...);
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output SEL;
    output SHIFT;
    output TDI;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCAN_VIRTEX5 (...);
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output SEL;
    output SHIFT;
    output TDI;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCAN_VIRTEX6 (...);
    parameter DISABLE_JTAG = "FALSE";
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCANE2 (...);
    parameter DISABLE_JTAG = "FALSE";
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

module DNA_PORT (...);
    parameter [56:0] SIM_DNA_VALUE = 57'h0;
    output DOUT;
    input CLK;
    input DIN;
    input READ;
    input SHIFT;
endmodule

module DNA_PORTE2 (...);
    parameter [95:0] SIM_DNA_VALUE = 96'h000000000000000000000000;
    output DOUT;
    input CLK;
    input DIN;
    input READ;
    input SHIFT;
endmodule

module FRAME_ECC_VIRTEX4 (...);
    output ERROR;
    output [11:0] SYNDROME;
    output SYNDROMEVALID;
endmodule

module FRAME_ECC_VIRTEX5 (...);
    output CRCERROR;
    output ECCERROR;
    output SYNDROMEVALID;
    output [11:0] SYNDROME;
endmodule

module FRAME_ECC_VIRTEX6 (...);
    parameter FARSRC = "EFAR";
    parameter FRAME_RBT_IN_FILENAME = "NONE";
    output CRCERROR;
    output ECCERROR;
    output ECCERRORSINGLE;
    output SYNDROMEVALID;
    output [12:0] SYNDROME;
    output [23:0] FAR;
    output [4:0] SYNBIT;
    output [6:0] SYNWORD;
endmodule

module FRAME_ECCE2 (...);
    parameter FARSRC = "EFAR";
    parameter FRAME_RBT_IN_FILENAME = "NONE";
    output CRCERROR;
    output ECCERROR;
    output ECCERRORSINGLE;
    output SYNDROMEVALID;
    output [12:0] SYNDROME;
    output [25:0] FAR;
    output [4:0] SYNBIT;
    output [6:0] SYNWORD;
endmodule

module FRAME_ECCE3 (...);
    output CRCERROR;
    output ECCERRORNOTSINGLE;
    output ECCERRORSINGLE;
    output ENDOFFRAME;
    output ENDOFSCAN;
    output [25:0] FAR;
    input [1:0] FARSEL;
    input ICAPBOTCLK;
    input ICAPTOPCLK;
endmodule

module USR_ACCESS_VIRTEX4 (...);
    output [31:0] DATA;
    output DATAVALID;
endmodule

module USR_ACCESS_VIRTEX5 (...);
    output CFGCLK;
    output [31:0] DATA;
    output DATAVALID;
endmodule

module USR_ACCESS_VIRTEX6 (...);
    output CFGCLK;
    output [31:0] DATA;
    output DATAVALID;
endmodule

module USR_ACCESSE2 (...);
    output CFGCLK;
    output DATAVALID;
    output [31:0] DATA;
endmodule

module POST_CRC_INTERNAL (...);
    output CRCERROR;
endmodule

(* keep *)
module SUSPEND_SYNC (...);
    output SREQ;
    input CLK;
    input SACK;
endmodule

(* keep *)
module KEY_CLEAR (...);
    input KEYCLEARB;
endmodule

(* keep *)
module MASTER_JTAG (...);
    output TDO;
    input TCK;
    input TDI;
    input TMS;
endmodule

(* keep *)
module SPI_ACCESS (...);
    parameter SIM_DELAY_TYPE = "SCALED";
    parameter SIM_DEVICE = "3S1400AN";
    parameter SIM_FACTORY_ID = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter SIM_MEM_FILE = "NONE";
    parameter SIM_USER_ID = 512'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    output MISO;
    input CLK;
    input CSB;
    input MOSI;
endmodule

module EFUSE_USR (...);
    parameter [31:0] SIM_EFUSE_VALUE = 32'h00000000;
    output [31:0] EFUSEUSR;
endmodule

module SYSMON (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0800;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter SIM_DEVICE = "VIRTEX5";
    parameter SIM_MONITOR_FILE = "design.txt";
    output BUSY;
    output DRDY;
    output EOC;
    output EOS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output OT;
    output [15:0] DO;
    output [2:0] ALM;
    output [4:0] CHANNEL;
    input CONVST;
    input CONVSTCLK;
    input DCLK;
    input DEN;
    input DWE;
    input RESET;
    input VN;
    input VP;
    input [15:0] DI;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input [6:0] DADDR;
endmodule

module XADC (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0800;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter [15:0] INIT_58 = 16'h0;
    parameter [15:0] INIT_59 = 16'h0;
    parameter [15:0] INIT_5A = 16'h0;
    parameter [15:0] INIT_5B = 16'h0;
    parameter [15:0] INIT_5C = 16'h0;
    parameter [15:0] INIT_5D = 16'h0;
    parameter [15:0] INIT_5E = 16'h0;
    parameter [15:0] INIT_5F = 16'h0;
    parameter IS_CONVSTCLK_INVERTED = 1'b0;
    parameter IS_DCLK_INVERTED = 1'b0;
    parameter SIM_DEVICE = "7SERIES";
    parameter SIM_MONITOR_FILE = "design.txt";
    output BUSY;
    output DRDY;
    output EOC;
    output EOS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output OT;
    output [15:0] DO;
    output [7:0] ALM;
    output [4:0] CHANNEL;
    output [4:0] MUXADDR;
    input CONVST;
    (* invertible_pin = "IS_CONVSTCLK_INVERTED" *)
    input CONVSTCLK;
    (* invertible_pin = "IS_DCLK_INVERTED" *)
    input DCLK;
    input DEN;
    input DWE;
    input RESET;
    input VN;
    input VP;
    input [15:0] DI;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input [6:0] DADDR;
endmodule

module SYSMONE1 (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter [15:0] INIT_58 = 16'h0;
    parameter [15:0] INIT_59 = 16'h0;
    parameter [15:0] INIT_5A = 16'h0;
    parameter [15:0] INIT_5B = 16'h0;
    parameter [15:0] INIT_5C = 16'h0;
    parameter [15:0] INIT_5D = 16'h0;
    parameter [15:0] INIT_5E = 16'h0;
    parameter [15:0] INIT_5F = 16'h0;
    parameter [15:0] INIT_60 = 16'h0;
    parameter [15:0] INIT_61 = 16'h0;
    parameter [15:0] INIT_62 = 16'h0;
    parameter [15:0] INIT_63 = 16'h0;
    parameter [15:0] INIT_64 = 16'h0;
    parameter [15:0] INIT_65 = 16'h0;
    parameter [15:0] INIT_66 = 16'h0;
    parameter [15:0] INIT_67 = 16'h0;
    parameter [15:0] INIT_68 = 16'h0;
    parameter [15:0] INIT_69 = 16'h0;
    parameter [15:0] INIT_6A = 16'h0;
    parameter [15:0] INIT_6B = 16'h0;
    parameter [15:0] INIT_6C = 16'h0;
    parameter [15:0] INIT_6D = 16'h0;
    parameter [15:0] INIT_6E = 16'h0;
    parameter [15:0] INIT_6F = 16'h0;
    parameter [15:0] INIT_70 = 16'h0;
    parameter [15:0] INIT_71 = 16'h0;
    parameter [15:0] INIT_72 = 16'h0;
    parameter [15:0] INIT_73 = 16'h0;
    parameter [15:0] INIT_74 = 16'h0;
    parameter [15:0] INIT_75 = 16'h0;
    parameter [15:0] INIT_76 = 16'h0;
    parameter [15:0] INIT_77 = 16'h0;
    parameter [15:0] INIT_78 = 16'h0;
    parameter [15:0] INIT_79 = 16'h0;
    parameter [15:0] INIT_7A = 16'h0;
    parameter [15:0] INIT_7B = 16'h0;
    parameter [15:0] INIT_7C = 16'h0;
    parameter [15:0] INIT_7D = 16'h0;
    parameter [15:0] INIT_7E = 16'h0;
    parameter [15:0] INIT_7F = 16'h0;
    parameter [0:0] IS_CONVSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DCLK_INVERTED = 1'b0;
    parameter SIM_MONITOR_FILE = "design.txt";
    parameter integer SYSMON_VUSER0_BANK = 0;
    parameter SYSMON_VUSER0_MONITOR = "NONE";
    parameter integer SYSMON_VUSER1_BANK = 0;
    parameter SYSMON_VUSER1_MONITOR = "NONE";
    parameter integer SYSMON_VUSER2_BANK = 0;
    parameter SYSMON_VUSER2_MONITOR = "NONE";
    parameter integer SYSMON_VUSER3_BANK = 0;
    parameter SYSMON_VUSER3_MONITOR = "NONE";
    output [15:0] ALM;
    output BUSY;
    output [5:0] CHANNEL;
    output [15:0] DO;
    output DRDY;
    output EOC;
    output EOS;
    output I2C_SCLK_TS;
    output I2C_SDA_TS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output [4:0] MUXADDR;
    output OT;
    input CONVST;
    (* invertible_pin = "IS_CONVSTCLK_INVERTED" *)
    input CONVSTCLK;
    input [7:0] DADDR;
    (* invertible_pin = "IS_DCLK_INVERTED" *)
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input I2C_SCLK;
    input I2C_SDA;
    input RESET;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input VN;
    input VP;
endmodule

module SYSMONE4 (...);
    parameter [15:0] COMMON_N_SOURCE = 16'hFFFF;
    parameter [15:0] INIT_40 = 16'h0000;
    parameter [15:0] INIT_41 = 16'h0000;
    parameter [15:0] INIT_42 = 16'h0000;
    parameter [15:0] INIT_43 = 16'h0000;
    parameter [15:0] INIT_44 = 16'h0000;
    parameter [15:0] INIT_45 = 16'h0000;
    parameter [15:0] INIT_46 = 16'h0000;
    parameter [15:0] INIT_47 = 16'h0000;
    parameter [15:0] INIT_48 = 16'h0000;
    parameter [15:0] INIT_49 = 16'h0000;
    parameter [15:0] INIT_4A = 16'h0000;
    parameter [15:0] INIT_4B = 16'h0000;
    parameter [15:0] INIT_4C = 16'h0000;
    parameter [15:0] INIT_4D = 16'h0000;
    parameter [15:0] INIT_4E = 16'h0000;
    parameter [15:0] INIT_4F = 16'h0000;
    parameter [15:0] INIT_50 = 16'h0000;
    parameter [15:0] INIT_51 = 16'h0000;
    parameter [15:0] INIT_52 = 16'h0000;
    parameter [15:0] INIT_53 = 16'h0000;
    parameter [15:0] INIT_54 = 16'h0000;
    parameter [15:0] INIT_55 = 16'h0000;
    parameter [15:0] INIT_56 = 16'h0000;
    parameter [15:0] INIT_57 = 16'h0000;
    parameter [15:0] INIT_58 = 16'h0000;
    parameter [15:0] INIT_59 = 16'h0000;
    parameter [15:0] INIT_5A = 16'h0000;
    parameter [15:0] INIT_5B = 16'h0000;
    parameter [15:0] INIT_5C = 16'h0000;
    parameter [15:0] INIT_5D = 16'h0000;
    parameter [15:0] INIT_5E = 16'h0000;
    parameter [15:0] INIT_5F = 16'h0000;
    parameter [15:0] INIT_60 = 16'h0000;
    parameter [15:0] INIT_61 = 16'h0000;
    parameter [15:0] INIT_62 = 16'h0000;
    parameter [15:0] INIT_63 = 16'h0000;
    parameter [15:0] INIT_64 = 16'h0000;
    parameter [15:0] INIT_65 = 16'h0000;
    parameter [15:0] INIT_66 = 16'h0000;
    parameter [15:0] INIT_67 = 16'h0000;
    parameter [15:0] INIT_68 = 16'h0000;
    parameter [15:0] INIT_69 = 16'h0000;
    parameter [15:0] INIT_6A = 16'h0000;
    parameter [15:0] INIT_6B = 16'h0000;
    parameter [15:0] INIT_6C = 16'h0000;
    parameter [15:0] INIT_6D = 16'h0000;
    parameter [15:0] INIT_6E = 16'h0000;
    parameter [15:0] INIT_6F = 16'h0000;
    parameter [15:0] INIT_70 = 16'h0000;
    parameter [15:0] INIT_71 = 16'h0000;
    parameter [15:0] INIT_72 = 16'h0000;
    parameter [15:0] INIT_73 = 16'h0000;
    parameter [15:0] INIT_74 = 16'h0000;
    parameter [15:0] INIT_75 = 16'h0000;
    parameter [15:0] INIT_76 = 16'h0000;
    parameter [15:0] INIT_77 = 16'h0000;
    parameter [15:0] INIT_78 = 16'h0000;
    parameter [15:0] INIT_79 = 16'h0000;
    parameter [15:0] INIT_7A = 16'h0000;
    parameter [15:0] INIT_7B = 16'h0000;
    parameter [15:0] INIT_7C = 16'h0000;
    parameter [15:0] INIT_7D = 16'h0000;
    parameter [15:0] INIT_7E = 16'h0000;
    parameter [15:0] INIT_7F = 16'h0000;
    parameter [0:0] IS_CONVSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DCLK_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MONITOR_FILE = "design.txt";
    parameter integer SYSMON_VUSER0_BANK = 0;
    parameter SYSMON_VUSER0_MONITOR = "NONE";
    parameter integer SYSMON_VUSER1_BANK = 0;
    parameter SYSMON_VUSER1_MONITOR = "NONE";
    parameter integer SYSMON_VUSER2_BANK = 0;
    parameter SYSMON_VUSER2_MONITOR = "NONE";
    parameter integer SYSMON_VUSER3_BANK = 0;
    parameter SYSMON_VUSER3_MONITOR = "NONE";
    output [15:0] ADC_DATA;
    output [15:0] ALM;
    output BUSY;
    output [5:0] CHANNEL;
    output [15:0] DO;
    output DRDY;
    output EOC;
    output EOS;
    output I2C_SCLK_TS;
    output I2C_SDA_TS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output [4:0] MUXADDR;
    output OT;
    output SMBALERT_TS;
    input CONVST;
    (* invertible_pin = "IS_CONVSTCLK_INVERTED" *)
    input CONVSTCLK;
    input [7:0] DADDR;
    (* invertible_pin = "IS_DCLK_INVERTED" *)
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input I2C_SCLK;
    input I2C_SDA;
    input RESET;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input VN;
    input VP;
endmodule

module GTPA1_DUAL (...);
    parameter AC_CAP_DIS_0 = "TRUE";
    parameter AC_CAP_DIS_1 = "TRUE";
    parameter integer ALIGN_COMMA_WORD_0 = 1;
    parameter integer ALIGN_COMMA_WORD_1 = 1;
    parameter integer CB2_INH_CC_PERIOD_0 = 8;
    parameter integer CB2_INH_CC_PERIOD_1 = 8;
    parameter [4:0] CDR_PH_ADJ_TIME_0 = 5'b01010;
    parameter [4:0] CDR_PH_ADJ_TIME_1 = 5'b01010;
    parameter integer CHAN_BOND_1_MAX_SKEW_0 = 7;
    parameter integer CHAN_BOND_1_MAX_SKEW_1 = 7;
    parameter integer CHAN_BOND_2_MAX_SKEW_0 = 1;
    parameter integer CHAN_BOND_2_MAX_SKEW_1 = 1;
    parameter CHAN_BOND_KEEP_ALIGN_0 = "FALSE";
    parameter CHAN_BOND_KEEP_ALIGN_1 = "FALSE";
    parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE_0 = "FALSE";
    parameter CHAN_BOND_SEQ_2_USE_1 = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN_0 = 1;
    parameter integer CHAN_BOND_SEQ_LEN_1 = 1;
    parameter integer CLK25_DIVIDER_0 = 4;
    parameter integer CLK25_DIVIDER_1 = 4;
    parameter CLKINDC_B_0 = "TRUE";
    parameter CLKINDC_B_1 = "TRUE";
    parameter CLKRCV_TRST_0 = "TRUE";
    parameter CLKRCV_TRST_1 = "TRUE";
    parameter CLK_CORRECT_USE_0 = "TRUE";
    parameter CLK_CORRECT_USE_1 = "TRUE";
    parameter integer CLK_COR_ADJ_LEN_0 = 1;
    parameter integer CLK_COR_ADJ_LEN_1 = 1;
    parameter integer CLK_COR_DET_LEN_0 = 1;
    parameter integer CLK_COR_DET_LEN_1 = 1;
    parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
    parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
    parameter integer CLK_COR_MAX_LAT_0 = 20;
    parameter integer CLK_COR_MAX_LAT_1 = 20;
    parameter integer CLK_COR_MIN_LAT_0 = 18;
    parameter integer CLK_COR_MIN_LAT_1 = 18;
    parameter CLK_COR_PRECEDENCE_0 = "TRUE";
    parameter CLK_COR_PRECEDENCE_1 = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT_0 = 0;
    parameter integer CLK_COR_REPEAT_WAIT_1 = 0;
    parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
    parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
    parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
    parameter CLK_OUT_GTP_SEL_0 = "REFCLKPLL0";
    parameter CLK_OUT_GTP_SEL_1 = "REFCLKPLL1";
    parameter [1:0] CM_TRIM_0 = 2'b00;
    parameter [1:0] CM_TRIM_1 = 2'b00;
    parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
    parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
    parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
    parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
    parameter DEC_MCOMMA_DETECT_0 = "TRUE";
    parameter DEC_MCOMMA_DETECT_1 = "TRUE";
    parameter DEC_PCOMMA_DETECT_0 = "TRUE";
    parameter DEC_PCOMMA_DETECT_1 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
    parameter GTP_CFG_PWRUP_0 = "TRUE";
    parameter GTP_CFG_PWRUP_1 = "TRUE";
    parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
    parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
    parameter MCOMMA_DETECT_0 = "TRUE";
    parameter MCOMMA_DETECT_1 = "TRUE";
    parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b110;
    parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b110;
    parameter integer OOB_CLK_DIVIDER_0 = 4;
    parameter integer OOB_CLK_DIVIDER_1 = 4;
    parameter PCI_EXPRESS_MODE_0 = "FALSE";
    parameter PCI_EXPRESS_MODE_1 = "FALSE";
    parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
    parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
    parameter PCOMMA_DETECT_0 = "TRUE";
    parameter PCOMMA_DETECT_1 = "TRUE";
    parameter [2:0] PLLLKDET_CFG_0 = 3'b101;
    parameter [2:0] PLLLKDET_CFG_1 = 3'b101;
    parameter [23:0] PLL_COM_CFG_0 = 24'h21680A;
    parameter [23:0] PLL_COM_CFG_1 = 24'h21680A;
    parameter [7:0] PLL_CP_CFG_0 = 8'h00;
    parameter [7:0] PLL_CP_CFG_1 = 8'h00;
    parameter integer PLL_DIVSEL_FB_0 = 5;
    parameter integer PLL_DIVSEL_FB_1 = 5;
    parameter integer PLL_DIVSEL_REF_0 = 2;
    parameter integer PLL_DIVSEL_REF_1 = 2;
    parameter integer PLL_RXDIVSEL_OUT_0 = 1;
    parameter integer PLL_RXDIVSEL_OUT_1 = 1;
    parameter PLL_SATA_0 = "FALSE";
    parameter PLL_SATA_1 = "FALSE";
    parameter PLL_SOURCE_0 = "PLL0";
    parameter PLL_SOURCE_1 = "PLL0";
    parameter integer PLL_TXDIVSEL_OUT_0 = 1;
    parameter integer PLL_TXDIVSEL_OUT_1 = 1;
    parameter [26:0] PMA_CDR_SCAN_0 = 27'h6404040;
    parameter [26:0] PMA_CDR_SCAN_1 = 27'h6404040;
    parameter [35:0] PMA_COM_CFG_EAST = 36'h000008000;
    parameter [35:0] PMA_COM_CFG_WEST = 36'h00000A000;
    parameter [6:0] PMA_RXSYNC_CFG_0 = 7'h00;
    parameter [6:0] PMA_RXSYNC_CFG_1 = 7'h00;
    parameter [24:0] PMA_RX_CFG_0 = 25'h05CE048;
    parameter [24:0] PMA_RX_CFG_1 = 25'h05CE048;
    parameter [19:0] PMA_TX_CFG_0 = 20'h00082;
    parameter [19:0] PMA_TX_CFG_1 = 20'h00082;
    parameter RCV_TERM_GND_0 = "FALSE";
    parameter RCV_TERM_GND_1 = "FALSE";
    parameter RCV_TERM_VTTRX_0 = "TRUE";
    parameter RCV_TERM_VTTRX_1 = "TRUE";
    parameter [7:0] RXEQ_CFG_0 = 8'b01111011;
    parameter [7:0] RXEQ_CFG_1 = 8'b01111011;
    parameter [0:0] RXPRBSERR_LOOPBACK_0 = 1'b0;
    parameter [0:0] RXPRBSERR_LOOPBACK_1 = 1'b0;
    parameter RX_BUFFER_USE_0 = "TRUE";
    parameter RX_BUFFER_USE_1 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
    parameter RX_EN_IDLE_HOLD_CDR_0 = "FALSE";
    parameter RX_EN_IDLE_HOLD_CDR_1 = "FALSE";
    parameter RX_EN_IDLE_RESET_BUF_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_BUF_1 = "TRUE";
    parameter RX_EN_IDLE_RESET_FR_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_FR_1 = "TRUE";
    parameter RX_EN_IDLE_RESET_PH_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_PH_1 = "TRUE";
    parameter RX_EN_MODE_RESET_BUF_0 = "TRUE";
    parameter RX_EN_MODE_RESET_BUF_1 = "TRUE";
    parameter [3:0] RX_IDLE_HI_CNT_0 = 4'b1000;
    parameter [3:0] RX_IDLE_HI_CNT_1 = 4'b1000;
    parameter [3:0] RX_IDLE_LO_CNT_0 = 4'b0000;
    parameter [3:0] RX_IDLE_LO_CNT_1 = 4'b0000;
    parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
    parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
    parameter integer RX_LOS_INVALID_INCR_0 = 1;
    parameter integer RX_LOS_INVALID_INCR_1 = 1;
    parameter integer RX_LOS_THRESHOLD_0 = 4;
    parameter integer RX_LOS_THRESHOLD_1 = 4;
    parameter RX_SLIDE_MODE_0 = "PCS";
    parameter RX_SLIDE_MODE_1 = "PCS";
    parameter RX_STATUS_FMT_0 = "PCIE";
    parameter RX_STATUS_FMT_1 = "PCIE";
    parameter RX_XCLK_SEL_0 = "RXREC";
    parameter RX_XCLK_SEL_1 = "RXREC";
    parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
    parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
    parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
    parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
    parameter integer SATA_MAX_BURST_0 = 7;
    parameter integer SATA_MAX_BURST_1 = 7;
    parameter integer SATA_MAX_INIT_0 = 22;
    parameter integer SATA_MAX_INIT_1 = 22;
    parameter integer SATA_MAX_WAKE_0 = 7;
    parameter integer SATA_MAX_WAKE_1 = 7;
    parameter integer SATA_MIN_BURST_0 = 4;
    parameter integer SATA_MIN_BURST_1 = 4;
    parameter integer SATA_MIN_INIT_0 = 12;
    parameter integer SATA_MIN_INIT_1 = 12;
    parameter integer SATA_MIN_WAKE_0 = 4;
    parameter integer SATA_MIN_WAKE_1 = 4;
    parameter integer SIM_GTPRESET_SPEEDUP = 0;
    parameter SIM_RECEIVER_DETECT_PASS = "FALSE";
    parameter [2:0] SIM_REFCLK0_SOURCE = 3'b000;
    parameter [2:0] SIM_REFCLK1_SOURCE = 3'b000;
    parameter SIM_TX_ELEC_IDLE_LEVEL = "X";
    parameter SIM_VERSION = "2.0";
    parameter [4:0] TERMINATION_CTRL_0 = 5'b10100;
    parameter [4:0] TERMINATION_CTRL_1 = 5'b10100;
    parameter TERMINATION_OVRD_0 = "FALSE";
    parameter TERMINATION_OVRD_1 = "FALSE";
    parameter [11:0] TRANS_TIME_FROM_P2_0 = 12'h03C;
    parameter [11:0] TRANS_TIME_FROM_P2_1 = 12'h03C;
    parameter [7:0] TRANS_TIME_NON_P2_0 = 8'h19;
    parameter [7:0] TRANS_TIME_NON_P2_1 = 8'h19;
    parameter [9:0] TRANS_TIME_TO_P2_0 = 10'h064;
    parameter [9:0] TRANS_TIME_TO_P2_1 = 10'h064;
    parameter [31:0] TST_ATTR_0 = 32'h00000000;
    parameter [31:0] TST_ATTR_1 = 32'h00000000;
    parameter [2:0] TXRX_INVERT_0 = 3'b011;
    parameter [2:0] TXRX_INVERT_1 = 3'b011;
    parameter TX_BUFFER_USE_0 = "FALSE";
    parameter TX_BUFFER_USE_1 = "FALSE";
    parameter [13:0] TX_DETECT_RX_CFG_0 = 14'h1832;
    parameter [13:0] TX_DETECT_RX_CFG_1 = 14'h1832;
    parameter [2:0] TX_IDLE_DELAY_0 = 3'b011;
    parameter [2:0] TX_IDLE_DELAY_1 = 3'b011;
    parameter [1:0] TX_TDCC_CFG_0 = 2'b00;
    parameter [1:0] TX_TDCC_CFG_1 = 2'b00;
    parameter TX_XCLK_SEL_0 = "TXUSR";
    parameter TX_XCLK_SEL_1 = "TXUSR";
    output DRDY;
    output PHYSTATUS0;
    output PHYSTATUS1;
    output PLLLKDET0;
    output PLLLKDET1;
    output REFCLKOUT0;
    output REFCLKOUT1;
    output REFCLKPLL0;
    output REFCLKPLL1;
    output RESETDONE0;
    output RESETDONE1;
    output RXBYTEISALIGNED0;
    output RXBYTEISALIGNED1;
    output RXBYTEREALIGN0;
    output RXBYTEREALIGN1;
    output RXCHANBONDSEQ0;
    output RXCHANBONDSEQ1;
    output RXCHANISALIGNED0;
    output RXCHANISALIGNED1;
    output RXCHANREALIGN0;
    output RXCHANREALIGN1;
    output RXCOMMADET0;
    output RXCOMMADET1;
    output RXELECIDLE0;
    output RXELECIDLE1;
    output RXPRBSERR0;
    output RXPRBSERR1;
    output RXRECCLK0;
    output RXRECCLK1;
    output RXVALID0;
    output RXVALID1;
    output TXN0;
    output TXN1;
    output TXOUTCLK0;
    output TXOUTCLK1;
    output TXP0;
    output TXP1;
    output [15:0] DRPDO;
    output [1:0] GTPCLKFBEAST;
    output [1:0] GTPCLKFBWEST;
    output [1:0] GTPCLKOUT0;
    output [1:0] GTPCLKOUT1;
    output [1:0] RXLOSSOFSYNC0;
    output [1:0] RXLOSSOFSYNC1;
    output [1:0] TXBUFSTATUS0;
    output [1:0] TXBUFSTATUS1;
    output [2:0] RXBUFSTATUS0;
    output [2:0] RXBUFSTATUS1;
    output [2:0] RXCHBONDO;
    output [2:0] RXCLKCORCNT0;
    output [2:0] RXCLKCORCNT1;
    output [2:0] RXSTATUS0;
    output [2:0] RXSTATUS1;
    output [31:0] RXDATA0;
    output [31:0] RXDATA1;
    output [3:0] RXCHARISCOMMA0;
    output [3:0] RXCHARISCOMMA1;
    output [3:0] RXCHARISK0;
    output [3:0] RXCHARISK1;
    output [3:0] RXDISPERR0;
    output [3:0] RXDISPERR1;
    output [3:0] RXNOTINTABLE0;
    output [3:0] RXNOTINTABLE1;
    output [3:0] RXRUNDISP0;
    output [3:0] RXRUNDISP1;
    output [3:0] TXKERR0;
    output [3:0] TXKERR1;
    output [3:0] TXRUNDISP0;
    output [3:0] TXRUNDISP1;
    output [4:0] RCALOUTEAST;
    output [4:0] RCALOUTWEST;
    output [4:0] TSTOUT0;
    output [4:0] TSTOUT1;
    input CLK00;
    input CLK01;
    input CLK10;
    input CLK11;
    input CLKINEAST0;
    input CLKINEAST1;
    input CLKINWEST0;
    input CLKINWEST1;
    input DCLK;
    input DEN;
    input DWE;
    input GATERXELECIDLE0;
    input GATERXELECIDLE1;
    input GCLK00;
    input GCLK01;
    input GCLK10;
    input GCLK11;
    input GTPRESET0;
    input GTPRESET1;
    input IGNORESIGDET0;
    input IGNORESIGDET1;
    input INTDATAWIDTH0;
    input INTDATAWIDTH1;
    input PLLCLK00;
    input PLLCLK01;
    input PLLCLK10;
    input PLLCLK11;
    input PLLLKDETEN0;
    input PLLLKDETEN1;
    input PLLPOWERDOWN0;
    input PLLPOWERDOWN1;
    input PRBSCNTRESET0;
    input PRBSCNTRESET1;
    input REFCLKPWRDNB0;
    input REFCLKPWRDNB1;
    input RXBUFRESET0;
    input RXBUFRESET1;
    input RXCDRRESET0;
    input RXCDRRESET1;
    input RXCHBONDMASTER0;
    input RXCHBONDMASTER1;
    input RXCHBONDSLAVE0;
    input RXCHBONDSLAVE1;
    input RXCOMMADETUSE0;
    input RXCOMMADETUSE1;
    input RXDEC8B10BUSE0;
    input RXDEC8B10BUSE1;
    input RXENCHANSYNC0;
    input RXENCHANSYNC1;
    input RXENMCOMMAALIGN0;
    input RXENMCOMMAALIGN1;
    input RXENPCOMMAALIGN0;
    input RXENPCOMMAALIGN1;
    input RXENPMAPHASEALIGN0;
    input RXENPMAPHASEALIGN1;
    input RXN0;
    input RXN1;
    input RXP0;
    input RXP1;
    input RXPMASETPHASE0;
    input RXPMASETPHASE1;
    input RXPOLARITY0;
    input RXPOLARITY1;
    input RXRESET0;
    input RXRESET1;
    input RXSLIDE0;
    input RXSLIDE1;
    input RXUSRCLK0;
    input RXUSRCLK1;
    input RXUSRCLK20;
    input RXUSRCLK21;
    input TSTCLK0;
    input TSTCLK1;
    input TXCOMSTART0;
    input TXCOMSTART1;
    input TXCOMTYPE0;
    input TXCOMTYPE1;
    input TXDETECTRX0;
    input TXDETECTRX1;
    input TXELECIDLE0;
    input TXELECIDLE1;
    input TXENC8B10BUSE0;
    input TXENC8B10BUSE1;
    input TXENPMAPHASEALIGN0;
    input TXENPMAPHASEALIGN1;
    input TXINHIBIT0;
    input TXINHIBIT1;
    input TXPDOWNASYNCH0;
    input TXPDOWNASYNCH1;
    input TXPMASETPHASE0;
    input TXPMASETPHASE1;
    input TXPOLARITY0;
    input TXPOLARITY1;
    input TXPRBSFORCEERR0;
    input TXPRBSFORCEERR1;
    input TXRESET0;
    input TXRESET1;
    input TXUSRCLK0;
    input TXUSRCLK1;
    input TXUSRCLK20;
    input TXUSRCLK21;
    input USRCODEERR0;
    input USRCODEERR1;
    input [11:0] TSTIN0;
    input [11:0] TSTIN1;
    input [15:0] DI;
    input [1:0] GTPCLKFBSEL0EAST;
    input [1:0] GTPCLKFBSEL0WEST;
    input [1:0] GTPCLKFBSEL1EAST;
    input [1:0] GTPCLKFBSEL1WEST;
    input [1:0] RXDATAWIDTH0;
    input [1:0] RXDATAWIDTH1;
    input [1:0] RXEQMIX0;
    input [1:0] RXEQMIX1;
    input [1:0] RXPOWERDOWN0;
    input [1:0] RXPOWERDOWN1;
    input [1:0] TXDATAWIDTH0;
    input [1:0] TXDATAWIDTH1;
    input [1:0] TXPOWERDOWN0;
    input [1:0] TXPOWERDOWN1;
    input [2:0] LOOPBACK0;
    input [2:0] LOOPBACK1;
    input [2:0] REFSELDYPLL0;
    input [2:0] REFSELDYPLL1;
    input [2:0] RXCHBONDI;
    input [2:0] RXENPRBSTST0;
    input [2:0] RXENPRBSTST1;
    input [2:0] TXBUFDIFFCTRL0;
    input [2:0] TXBUFDIFFCTRL1;
    input [2:0] TXENPRBSTST0;
    input [2:0] TXENPRBSTST1;
    input [2:0] TXPREEMPHASIS0;
    input [2:0] TXPREEMPHASIS1;
    input [31:0] TXDATA0;
    input [31:0] TXDATA1;
    input [3:0] TXBYPASS8B10B0;
    input [3:0] TXBYPASS8B10B1;
    input [3:0] TXCHARDISPMODE0;
    input [3:0] TXCHARDISPMODE1;
    input [3:0] TXCHARDISPVAL0;
    input [3:0] TXCHARDISPVAL1;
    input [3:0] TXCHARISK0;
    input [3:0] TXCHARISK1;
    input [3:0] TXDIFFCTRL0;
    input [3:0] TXDIFFCTRL1;
    input [4:0] RCALINEAST;
    input [4:0] RCALINWEST;
    input [7:0] DADDR;
    input [7:0] GTPTEST0;
    input [7:0] GTPTEST1;
endmodule

module GT11_CUSTOM (...);
    parameter ALIGN_COMMA_WORD = 1;
    parameter BANDGAPSEL = "FALSE";
    parameter BIASRESSEL = "TRUE";
    parameter CCCB_ARBITRATOR_DISABLE = "FALSE";
    parameter CHAN_BOND_LIMIT = 16;
    parameter CHAN_BOND_MODE = "NONE";
    parameter CHAN_BOND_ONE_SHOT = "FALSE";
    parameter CHAN_BOND_SEQ_1_1 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_2 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_3 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_4 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_MASK = 4'b0000;
    parameter CHAN_BOND_SEQ_2_1 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_2 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_3 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_4 = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_MASK = 4'b0000;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_8B10B_DE = "FALSE";
    parameter CLK_COR_MAX_LAT = 36;
    parameter CLK_COR_MIN_LAT = 28;
    parameter CLK_COR_SEQ_1_1 = 11'b00000000000;
    parameter CLK_COR_SEQ_1_2 = 11'b00000000000;
    parameter CLK_COR_SEQ_1_3 = 11'b00000000000;
    parameter CLK_COR_SEQ_1_4 = 11'b00000000000;
    parameter CLK_COR_SEQ_1_MASK = 4'b0000;
    parameter CLK_COR_SEQ_2_1 = 11'b00000000000;
    parameter CLK_COR_SEQ_2_2 = 11'b00000000000;
    parameter CLK_COR_SEQ_2_3 = 11'b00000000000;
    parameter CLK_COR_SEQ_2_4 = 11'b00000000000;
    parameter CLK_COR_SEQ_2_MASK = 4'b0000;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter CLK_COR_SEQ_DROP = "FALSE";
    parameter CLK_COR_SEQ_LEN = 1;
    parameter COMMA32 = "FALSE";
    parameter COMMA_10B_MASK = 10'h3FF;
    parameter CYCLE_LIMIT_SEL = 2'b00;
    parameter DCDR_FILTER = 3'b010;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter DIGRX_FWDCLK = 2'b00;
    parameter DIGRX_SYNC_MODE = "FALSE";
    parameter ENABLE_DCDR = "FALSE";
    parameter FDET_HYS_CAL = 3'b110;
    parameter FDET_HYS_SEL = 3'b110;
    parameter FDET_LCK_CAL = 3'b101;
    parameter FDET_LCK_SEL = 3'b101;
    parameter GT11_MODE = "SINGLE";
    parameter IREFBIASMODE = 2'b11;
    parameter LOOPCAL_WAIT = 2'b00;
    parameter MCOMMA_32B_VALUE = 32'h000000F6;
    parameter MCOMMA_DETECT = "TRUE";
    parameter OPPOSITE_SELECT = "FALSE";
    parameter PCOMMA_32B_VALUE = 32'hF6F62828;
    parameter PCOMMA_DETECT = "TRUE";
    parameter PCS_BIT_SLIP = "FALSE";
    parameter PMACLKENABLE = "TRUE";
    parameter PMACOREPWRENABLE = "TRUE";
    parameter PMAIREFTRIM = 4'b0111;
    parameter PMAVBGCTRL = 5'b00000;
    parameter PMAVREFTRIM = 4'b0111;
    parameter PMA_BIT_SLIP = "FALSE";
    parameter REPEATER = "FALSE";
    parameter RXACTST = "FALSE";
    parameter RXAFEEQ = 9'b000000000;
    parameter RXAFEPD = "FALSE";
    parameter RXAFETST = "FALSE";
    parameter RXAPD = "FALSE";
    parameter RXASYNCDIVIDE = 2'b11;
    parameter RXBY_32 = "TRUE";
    parameter RXCDRLOS = 6'b000000;
    parameter RXCLK0_FORCE_PMACLK = "FALSE";
    parameter RXCLKMODE = 6'b110001;
    parameter RXCMADJ = 2'b10;
    parameter RXCPSEL = "TRUE";
    parameter RXCPTST = "FALSE";
    parameter RXCRCCLOCKDOUBLE = "FALSE";
    parameter RXCRCENABLE = "FALSE";
    parameter RXCRCINITVAL = 32'h00000000;
    parameter RXCRCINVERTGEN = "FALSE";
    parameter RXCRCSAMECLOCK = "FALSE";
    parameter RXCTRL1 = 10'h200;
    parameter RXCYCLE_LIMIT_SEL = 2'b00;
    parameter RXDATA_SEL = 2'b00;
    parameter RXDCCOUPLE = "FALSE";
    parameter RXDIGRESET = "FALSE";
    parameter RXDIGRX = "FALSE";
    parameter RXEQ = 64'h4000000000000000;
    parameter RXFDCAL_CLOCK_DIVIDE = "NONE";
    parameter RXFDET_HYS_CAL = 3'b110;
    parameter RXFDET_HYS_SEL = 3'b110;
    parameter RXFDET_LCK_CAL = 3'b101;
    parameter RXFDET_LCK_SEL = 3'b101;
    parameter RXFECONTROL1 = 2'b00;
    parameter RXFECONTROL2 = 3'b000;
    parameter RXFETUNE = 2'b01;
    parameter RXLB = "FALSE";
    parameter RXLKADJ = 5'b00000;
    parameter RXLKAPD = "FALSE";
    parameter RXLOOPCAL_WAIT = 2'b00;
    parameter RXLOOPFILT = 4'b0111;
    parameter RXOUTDIV2SEL = 1;
    parameter RXPD = "FALSE";
    parameter RXPDDTST = "FALSE";
    parameter RXPLLNDIVSEL = 8;
    parameter RXPMACLKSEL = "REFCLK1";
    parameter RXRCPADJ = 3'b011;
    parameter RXRCPPD = "FALSE";
    parameter RXRECCLK1_USE_SYNC = "FALSE";
    parameter RXRIBADJ = 2'b11;
    parameter RXRPDPD = "FALSE";
    parameter RXRSDPD = "FALSE";
    parameter RXSLOWDOWN_CAL = 2'b00;
    parameter RXUSRDIVISOR = 1;
    parameter RXVCODAC_INIT = 10'b1010000000;
    parameter RXVCO_CTRL_ENABLE = "TRUE";
    parameter RX_BUFFER_USE = "TRUE";
    parameter RX_CLOCK_DIVIDER = 2'b00;
    parameter RX_LOS_INVALID_INCR = 1;
    parameter RX_LOS_THRESHOLD = 4;
    parameter SAMPLE_8X = "FALSE";
    parameter SH_CNT_MAX = 64;
    parameter SH_INVALID_CNT_MAX = 16;
    parameter SLOWDOWN_CAL = 2'b00;
    parameter TXABPMACLKSEL = "REFCLK1";
    parameter TXAPD = "FALSE";
    parameter TXAREFBIASSEL = "FALSE";
    parameter TXASYNCDIVIDE = 2'b11;
    parameter TXCLK0_FORCE_PMACLK = "FALSE";
    parameter TXCLKMODE = 4'b1001;
    parameter TXCPSEL = "TRUE";
    parameter TXCRCCLOCKDOUBLE = "FALSE";
    parameter TXCRCENABLE = "FALSE";
    parameter TXCRCINITVAL = 32'h00000000;
    parameter TXCRCINVERTGEN = "FALSE";
    parameter TXCRCSAMECLOCK = "FALSE";
    parameter TXCTRL1 = 10'h200;
    parameter TXDATA_SEL = 2'b00;
    parameter TXDAT_PRDRV_DAC = 3'b111;
    parameter TXDAT_TAP_DAC = 5'b10110;
    parameter TXDIGPD = "FALSE";
    parameter TXFDCAL_CLOCK_DIVIDE = "NONE";
    parameter TXHIGHSIGNALEN = "TRUE";
    parameter TXLOOPFILT = 4'b0111;
    parameter TXLVLSHFTPD = "FALSE";
    parameter TXOUTCLK1_USE_SYNC = "FALSE";
    parameter TXOUTDIV2SEL = 1;
    parameter TXPD = "FALSE";
    parameter TXPHASESEL = "FALSE";
    parameter TXPLLNDIVSEL = 8;
    parameter TXPOST_PRDRV_DAC = 3'b111;
    parameter TXPOST_TAP_DAC = 5'b01110;
    parameter TXPOST_TAP_PD = "TRUE";
    parameter TXPRE_PRDRV_DAC = 3'b111;
    parameter TXPRE_TAP_DAC = 5'b00000;
    parameter TXPRE_TAP_PD = "TRUE";
    parameter TXSLEWRATE = "FALSE";
    parameter TXTERMTRIM = 4'b1100;
    parameter TX_BUFFER_USE = "TRUE";
    parameter TX_CLOCK_DIVIDER = 2'b00;
    parameter VCODAC_INIT = 10'b1010000000;
    parameter VCO_CTRL_ENABLE = "TRUE";
    parameter VREFBIASMODE = 2'b11;
    output DRDY;
    output RXBUFERR;
    output RXCALFAIL;
    output RXCOMMADET;
    output RXCYCLELIMIT;
    output RXLOCK;
    output RXMCLK;
    output RXPCSHCLKOUT;
    output RXREALIGN;
    output RXRECCLK1;
    output RXRECCLK2;
    output RXSIGDET;
    output TX1N;
    output TX1P;
    output TXBUFERR;
    output TXCALFAIL;
    output TXCYCLELIMIT;
    output TXLOCK;
    output TXOUTCLK1;
    output TXOUTCLK2;
    output TXPCSHCLKOUT;
    output [15:0] DO;
    output [1:0] RXLOSSOFSYNC;
    output [31:0] RXCRCOUT;
    output [31:0] TXCRCOUT;
    output [4:0] CHBONDO;
    output [5:0] RXSTATUS;
    output [63:0] RXDATA;
    output [7:0] RXCHARISCOMMA;
    output [7:0] RXCHARISK;
    output [7:0] RXDISPERR;
    output [7:0] RXNOTINTABLE;
    output [7:0] RXRUNDISP;
    output [7:0] TXKERR;
    output [7:0] TXRUNDISP;
    input DCLK;
    input DEN;
    input DWE;
    input ENCHANSYNC;
    input ENMCOMMAALIGN;
    input ENPCOMMAALIGN;
    input GREFCLK;
    input POWERDOWN;
    input REFCLK1;
    input REFCLK2;
    input RX1N;
    input RX1P;
    input RXBLOCKSYNC64B66BUSE;
    input RXCLKSTABLE;
    input RXCOMMADETUSE;
    input RXCRCCLK;
    input RXCRCDATAVALID;
    input RXCRCINIT;
    input RXCRCINTCLK;
    input RXCRCPD;
    input RXCRCRESET;
    input RXDEC64B66BUSE;
    input RXDEC8B10BUSE;
    input RXDESCRAM64B66BUSE;
    input RXIGNOREBTF;
    input RXPMARESET;
    input RXPOLARITY;
    input RXRESET;
    input RXSLIDE;
    input RXSYNC;
    input RXUSRCLK2;
    input RXUSRCLK;
    input TXCLKSTABLE;
    input TXCRCCLK;
    input TXCRCDATAVALID;
    input TXCRCINIT;
    input TXCRCINTCLK;
    input TXCRCPD;
    input TXCRCRESET;
    input TXENC64B66BUSE;
    input TXENC8B10BUSE;
    input TXENOOB;
    input TXGEARBOX64B66BUSE;
    input TXINHIBIT;
    input TXPMARESET;
    input TXPOLARITY;
    input TXRESET;
    input TXSCRAM64B66BUSE;
    input TXSYNC;
    input TXUSRCLK2;
    input TXUSRCLK;
    input [15:0] DI;
    input [1:0] LOOPBACK;
    input [1:0] RXDATAWIDTH;
    input [1:0] RXINTDATAWIDTH;
    input [1:0] TXDATAWIDTH;
    input [1:0] TXINTDATAWIDTH;
    input [2:0] RXCRCDATAWIDTH;
    input [2:0] TXCRCDATAWIDTH;
    input [4:0] CHBONDI;
    input [63:0] RXCRCIN;
    input [63:0] TXCRCIN;
    input [63:0] TXDATA;
    input [7:0] DADDR;
    input [7:0] TXBYPASS8B10B;
    input [7:0] TXCHARDISPMODE;
    input [7:0] TXCHARDISPVAL;
    input [7:0] TXCHARISK;
endmodule

module GT11_DUAL (...);
    parameter ALIGN_COMMA_WORD_A = 1;
    parameter ALIGN_COMMA_WORD_B = 1;
    parameter BANDGAPSEL_A = "FALSE";
    parameter BANDGAPSEL_B = "FALSE";
    parameter BIASRESSEL_A = "TRUE";
    parameter BIASRESSEL_B = "TRUE";
    parameter CCCB_ARBITRATOR_DISABLE_A = "FALSE";
    parameter CCCB_ARBITRATOR_DISABLE_B = "FALSE";
    parameter CHAN_BOND_LIMIT_A = 16;
    parameter CHAN_BOND_LIMIT_B = 16;
    parameter CHAN_BOND_MODE_A = "NONE";
    parameter CHAN_BOND_MODE_B = "NONE";
    parameter CHAN_BOND_ONE_SHOT_A = "FALSE";
    parameter CHAN_BOND_ONE_SHOT_B = "FALSE";
    parameter CHAN_BOND_SEQ_1_1_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_1_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_2_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_2_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_3_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_3_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_4_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_4_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_1_MASK_A = 4'b0000;
    parameter CHAN_BOND_SEQ_1_MASK_B = 4'b0000;
    parameter CHAN_BOND_SEQ_2_1_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_1_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_2_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_2_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_3_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_3_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_4_A = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_4_B = 11'b00000000000;
    parameter CHAN_BOND_SEQ_2_MASK_A = 4'b0000;
    parameter CHAN_BOND_SEQ_2_MASK_B = 4'b0000;
    parameter CHAN_BOND_SEQ_2_USE_A = "FALSE";
    parameter CHAN_BOND_SEQ_2_USE_B = "FALSE";
    parameter CHAN_BOND_SEQ_LEN_A = 1;
    parameter CHAN_BOND_SEQ_LEN_B = 1;
    parameter CLK_CORRECT_USE_A = "TRUE";
    parameter CLK_CORRECT_USE_B = "TRUE";
    parameter CLK_COR_8B10B_DE_A = "FALSE";
    parameter CLK_COR_8B10B_DE_B = "FALSE";
    parameter CLK_COR_MAX_LAT_A = 36;
    parameter CLK_COR_MAX_LAT_B = 36;
    parameter CLK_COR_MIN_LAT_A = 28;
    parameter CLK_COR_MIN_LAT_B = 28;
    parameter CLK_COR_SEQ_1_1_A = 11'b00000000000;
    parameter CLK_COR_SEQ_1_1_B = 11'b00000000000;
    parameter CLK_COR_SEQ_1_2_A = 11'b00000000000;
    parameter CLK_COR_SEQ_1_2_B = 11'b00000000000;
    parameter CLK_COR_SEQ_1_3_A = 11'b00000000000;
    parameter CLK_COR_SEQ_1_3_B = 11'b00000000000;
    parameter CLK_COR_SEQ_1_4_A = 11'b00000000000;
    parameter CLK_COR_SEQ_1_4_B = 11'b00000000000;
    parameter CLK_COR_SEQ_1_MASK_A = 4'b0000;
    parameter CLK_COR_SEQ_1_MASK_B = 4'b0000;
    parameter CLK_COR_SEQ_2_1_A = 11'b00000000000;
    parameter CLK_COR_SEQ_2_1_B = 11'b00000000000;
    parameter CLK_COR_SEQ_2_2_A = 11'b00000000000;
    parameter CLK_COR_SEQ_2_2_B = 11'b00000000000;
    parameter CLK_COR_SEQ_2_3_A = 11'b00000000000;
    parameter CLK_COR_SEQ_2_3_B = 11'b00000000000;
    parameter CLK_COR_SEQ_2_4_A = 11'b00000000000;
    parameter CLK_COR_SEQ_2_4_B = 11'b00000000000;
    parameter CLK_COR_SEQ_2_MASK_A = 4'b0000;
    parameter CLK_COR_SEQ_2_MASK_B = 4'b0000;
    parameter CLK_COR_SEQ_2_USE_A = "FALSE";
    parameter CLK_COR_SEQ_2_USE_B = "FALSE";
    parameter CLK_COR_SEQ_DROP_A = "FALSE";
    parameter CLK_COR_SEQ_DROP_B = "FALSE";
    parameter CLK_COR_SEQ_LEN_A = 1;
    parameter CLK_COR_SEQ_LEN_B = 1;
    parameter COMMA32_A = "FALSE";
    parameter COMMA32_B = "FALSE";
    parameter COMMA_10B_MASK_A = 10'h3FF;
    parameter COMMA_10B_MASK_B = 10'h3FF;
    parameter CYCLE_LIMIT_SEL_A = 2'b00;
    parameter CYCLE_LIMIT_SEL_B = 2'b00;
    parameter DCDR_FILTER_A = 3'b010;
    parameter DCDR_FILTER_B = 3'b010;
    parameter DEC_MCOMMA_DETECT_A = "TRUE";
    parameter DEC_MCOMMA_DETECT_B = "TRUE";
    parameter DEC_PCOMMA_DETECT_A = "TRUE";
    parameter DEC_PCOMMA_DETECT_B = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_A = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_B = "TRUE";
    parameter DIGRX_FWDCLK_A = 2'b00;
    parameter DIGRX_FWDCLK_B = 2'b00;
    parameter DIGRX_SYNC_MODE_A = "FALSE";
    parameter DIGRX_SYNC_MODE_B = "FALSE";
    parameter ENABLE_DCDR_A = "FALSE";
    parameter ENABLE_DCDR_B = "FALSE";
    parameter FDET_HYS_CAL_A = 3'b110;
    parameter FDET_HYS_CAL_B = 3'b110;
    parameter FDET_HYS_SEL_A = 3'b110;
    parameter FDET_HYS_SEL_B = 3'b110;
    parameter FDET_LCK_CAL_A = 3'b101;
    parameter FDET_LCK_CAL_B = 3'b101;
    parameter FDET_LCK_SEL_A = 3'b101;
    parameter FDET_LCK_SEL_B = 3'b101;
    parameter IREFBIASMODE_A = 2'b11;
    parameter IREFBIASMODE_B = 2'b11;
    parameter LOOPCAL_WAIT_A = 2'b00;
    parameter LOOPCAL_WAIT_B = 2'b00;
    parameter MCOMMA_32B_VALUE_A = 32'hA1A1A2A2;
    parameter MCOMMA_32B_VALUE_B = 32'hA1A1A2A2;
    parameter MCOMMA_DETECT_A = "TRUE";
    parameter MCOMMA_DETECT_B = "TRUE";
    parameter OPPOSITE_SELECT_A = "FALSE";
    parameter OPPOSITE_SELECT_B = "FALSE";
    parameter PCOMMA_32B_VALUE_A = 32'hA1A1A2A2;
    parameter PCOMMA_32B_VALUE_B = 32'hA1A1A2A2;
    parameter PCOMMA_DETECT_A = "TRUE";
    parameter PCOMMA_DETECT_B = "TRUE";
    parameter PCS_BIT_SLIP_A = "FALSE";
    parameter PCS_BIT_SLIP_B = "FALSE";
    parameter PMACLKENABLE_A = "TRUE";
    parameter PMACLKENABLE_B = "TRUE";
    parameter PMACOREPWRENABLE_A = "TRUE";
    parameter PMACOREPWRENABLE_B = "TRUE";
    parameter PMAIREFTRIM_A = 4'b0111;
    parameter PMAIREFTRIM_B = 4'b0111;
    parameter PMAVBGCTRL_A = 5'b00000;
    parameter PMAVBGCTRL_B = 5'b00000;
    parameter PMAVREFTRIM_A = 4'b0111;
    parameter PMAVREFTRIM_B = 4'b0111;
    parameter PMA_BIT_SLIP_A = "FALSE";
    parameter PMA_BIT_SLIP_B = "FALSE";
    parameter POWER_ENABLE_A = "TRUE";
    parameter POWER_ENABLE_B = "TRUE";
    parameter REPEATER_A = "FALSE";
    parameter REPEATER_B = "FALSE";
    parameter RXACTST_A = "FALSE";
    parameter RXACTST_B = "FALSE";
    parameter RXAFEEQ_A = 9'b000000000;
    parameter RXAFEEQ_B = 9'b000000000;
    parameter RXAFEPD_A = "FALSE";
    parameter RXAFEPD_B = "FALSE";
    parameter RXAFETST_A = "FALSE";
    parameter RXAFETST_B = "FALSE";
    parameter RXAPD_A = "FALSE";
    parameter RXAPD_B = "FALSE";
    parameter RXASYNCDIVIDE_A = 2'b00;
    parameter RXASYNCDIVIDE_B = 2'b00;
    parameter RXBY_32_A = "TRUE";
    parameter RXBY_32_B = "TRUE";
    parameter RXCDRLOS_A = 6'b000000;
    parameter RXCDRLOS_B = 6'b000000;
    parameter RXCLK0_FORCE_PMACLK_A = "FALSE";
    parameter RXCLK0_FORCE_PMACLK_B = "FALSE";
    parameter RXCLKMODE_A = 6'b110001;
    parameter RXCLKMODE_B = 6'b110001;
    parameter RXCMADJ_A = 2'b10;
    parameter RXCMADJ_B = 2'b10;
    parameter RXCPSEL_A = "TRUE";
    parameter RXCPSEL_B = "TRUE";
    parameter RXCPTST_A = "FALSE";
    parameter RXCPTST_B = "FALSE";
    parameter RXCRCCLOCKDOUBLE_A = "FALSE";
    parameter RXCRCCLOCKDOUBLE_B = "FALSE";
    parameter RXCRCENABLE_A = "FALSE";
    parameter RXCRCENABLE_B = "FALSE";
    parameter RXCRCINITVAL_A = 32'h00000000;
    parameter RXCRCINITVAL_B = 32'h00000000;
    parameter RXCRCINVERTGEN_A = "FALSE";
    parameter RXCRCINVERTGEN_B = "FALSE";
    parameter RXCRCSAMECLOCK_A = "FALSE";
    parameter RXCRCSAMECLOCK_B = "FALSE";
    parameter RXCTRL1_A = 10'h006;
    parameter RXCTRL1_B = 10'h006;
    parameter RXCYCLE_LIMIT_SEL_A = 2'b00;
    parameter RXCYCLE_LIMIT_SEL_B = 2'b00;
    parameter RXDATA_SEL_A = 2'b00;
    parameter RXDATA_SEL_B = 2'b00;
    parameter RXDCCOUPLE_A = "FALSE";
    parameter RXDCCOUPLE_B = "FALSE";
    parameter RXDIGRESET_A = "FALSE";
    parameter RXDIGRESET_B = "FALSE";
    parameter RXDIGRX_A = "FALSE";
    parameter RXDIGRX_B = "FALSE";
    parameter RXEQ_A = 64'h4000000000000000;
    parameter RXEQ_B = 64'h4000000000000000;
    parameter RXFDCAL_CLOCK_DIVIDE_A = "NONE";
    parameter RXFDCAL_CLOCK_DIVIDE_B = "NONE";
    parameter RXFDET_HYS_CAL_A = 3'b110;
    parameter RXFDET_HYS_CAL_B = 3'b110;
    parameter RXFDET_HYS_SEL_A = 3'b110;
    parameter RXFDET_HYS_SEL_B = 3'b110;
    parameter RXFDET_LCK_CAL_A = 3'b101;
    parameter RXFDET_LCK_CAL_B = 3'b101;
    parameter RXFDET_LCK_SEL_A = 3'b101;
    parameter RXFDET_LCK_SEL_B = 3'b101;
    parameter RXFECONTROL1_A = 2'b00;
    parameter RXFECONTROL1_B = 2'b00;
    parameter RXFECONTROL2_A = 3'b000;
    parameter RXFECONTROL2_B = 3'b000;
    parameter RXFETUNE_A = 2'b01;
    parameter RXFETUNE_B = 2'b01;
    parameter RXLB_A = "FALSE";
    parameter RXLB_B = "FALSE";
    parameter RXLKADJ_A = 5'b00000;
    parameter RXLKADJ_B = 5'b00000;
    parameter RXLKAPD_A = "FALSE";
    parameter RXLKAPD_B = "FALSE";
    parameter RXLOOPCAL_WAIT_A = 2'b00;
    parameter RXLOOPCAL_WAIT_B = 2'b00;
    parameter RXLOOPFILT_A = 4'b0111;
    parameter RXLOOPFILT_B = 4'b0111;
    parameter RXOUTDIV2SEL_A = 1;
    parameter RXOUTDIV2SEL_B = 1;
    parameter RXPDDTST_A = "FALSE";
    parameter RXPDDTST_B = "FALSE";
    parameter RXPD_A = "FALSE";
    parameter RXPD_B = "FALSE";
    parameter RXPLLNDIVSEL_A = 8;
    parameter RXPLLNDIVSEL_B = 8;
    parameter RXPMACLKSEL_A = "REFCLK1";
    parameter RXPMACLKSEL_B = "REFCLK1";
    parameter RXRCPADJ_A = 3'b011;
    parameter RXRCPADJ_B = 3'b011;
    parameter RXRCPPD_A = "FALSE";
    parameter RXRCPPD_B = "FALSE";
    parameter RXRECCLK1_USE_SYNC_A = "FALSE";
    parameter RXRECCLK1_USE_SYNC_B = "FALSE";
    parameter RXRIBADJ_A = 2'b11;
    parameter RXRIBADJ_B = 2'b11;
    parameter RXRPDPD_A = "FALSE";
    parameter RXRPDPD_B = "FALSE";
    parameter RXRSDPD_A = "FALSE";
    parameter RXRSDPD_B = "FALSE";
    parameter RXSLOWDOWN_CAL_A = 2'b00;
    parameter RXSLOWDOWN_CAL_B = 2'b00;
    parameter RXUSRDIVISOR_A = 1;
    parameter RXUSRDIVISOR_B = 1;
    parameter RXVCODAC_INIT_A = 10'b1010000000;
    parameter RXVCODAC_INIT_B = 10'b1010000000;
    parameter RXVCO_CTRL_ENABLE_A = "TRUE";
    parameter RXVCO_CTRL_ENABLE_B = "TRUE";
    parameter RX_BUFFER_USE_A = "TRUE";
    parameter RX_BUFFER_USE_B = "TRUE";
    parameter RX_CLOCK_DIVIDER_A = 2'b00;
    parameter RX_CLOCK_DIVIDER_B = 2'b00;
    parameter RX_LOS_INVALID_INCR_A = 1;
    parameter RX_LOS_INVALID_INCR_B = 1;
    parameter RX_LOS_THRESHOLD_A = 4;
    parameter RX_LOS_THRESHOLD_B = 4;
    parameter SAMPLE_8X_A = "FALSE";
    parameter SAMPLE_8X_B = "FALSE";
    parameter SH_CNT_MAX_A = 64;
    parameter SH_CNT_MAX_B = 64;
    parameter SH_INVALID_CNT_MAX_A = 16;
    parameter SH_INVALID_CNT_MAX_B = 16;
    parameter SLOWDOWN_CAL_A = 2'b00;
    parameter SLOWDOWN_CAL_B = 2'b00;
    parameter TXABPMACLKSEL_A = "REFCLK1";
    parameter TXABPMACLKSEL_B = "REFCLK1";
    parameter TXAPD_A = "FALSE";
    parameter TXAPD_B = "FALSE";
    parameter TXAREFBIASSEL_A = "FALSE";
    parameter TXAREFBIASSEL_B = "FALSE";
    parameter TXASYNCDIVIDE_A = 2'b00;
    parameter TXASYNCDIVIDE_B = 2'b00;
    parameter TXCLK0_FORCE_PMACLK_A = "FALSE";
    parameter TXCLK0_FORCE_PMACLK_B = "FALSE";
    parameter TXCLKMODE_A = 4'b1001;
    parameter TXCLKMODE_B = 4'b1001;
    parameter TXCPSEL_A = "TRUE";
    parameter TXCPSEL_B = "TRUE";
    parameter TXCRCCLOCKDOUBLE_A = "FALSE";
    parameter TXCRCCLOCKDOUBLE_B = "FALSE";
    parameter TXCRCENABLE_A = "FALSE";
    parameter TXCRCENABLE_B = "FALSE";
    parameter TXCRCINITVAL_A = 32'h00000000;
    parameter TXCRCINITVAL_B = 32'h00000000;
    parameter TXCRCINVERTGEN_A = "FALSE";
    parameter TXCRCINVERTGEN_B = "FALSE";
    parameter TXCRCSAMECLOCK_A = "FALSE";
    parameter TXCRCSAMECLOCK_B = "FALSE";
    parameter TXCTRL1_A = 10'h006;
    parameter TXCTRL1_B = 10'h006;
    parameter TXDATA_SEL_A = 2'b00;
    parameter TXDATA_SEL_B = 2'b00;
    parameter TXDAT_PRDRV_DAC_A = 3'b111;
    parameter TXDAT_PRDRV_DAC_B = 3'b111;
    parameter TXDAT_TAP_DAC_A = 5'b10110;
    parameter TXDAT_TAP_DAC_B = 5'b10110;
    parameter TXDIGPD_A = "FALSE";
    parameter TXDIGPD_B = "FALSE";
    parameter TXFDCAL_CLOCK_DIVIDE_A = "NONE";
    parameter TXFDCAL_CLOCK_DIVIDE_B = "NONE";
    parameter TXHIGHSIGNALEN_A = "TRUE";
    parameter TXHIGHSIGNALEN_B = "TRUE";
    parameter TXLOOPFILT_A = 4'b0111;
    parameter TXLOOPFILT_B = 4'b0111;
    parameter TXLVLSHFTPD_A = "FALSE";
    parameter TXLVLSHFTPD_B = "FALSE";
    parameter TXOUTCLK1_USE_SYNC_A = "FALSE";
    parameter TXOUTCLK1_USE_SYNC_B = "FALSE";
    parameter TXOUTDIV2SEL_A = 1;
    parameter TXOUTDIV2SEL_B = 1;
    parameter TXPD_A = "FALSE";
    parameter TXPD_B = "FALSE";
    parameter TXPHASESEL_A = "FALSE";
    parameter TXPHASESEL_B = "FALSE";
    parameter TXPLLNDIVSEL_A = 8;
    parameter TXPLLNDIVSEL_B = 8;
    parameter TXPOST_PRDRV_DAC_A = 3'b111;
    parameter TXPOST_PRDRV_DAC_B = 3'b111;
    parameter TXPOST_TAP_DAC_A = 5'b01110;
    parameter TXPOST_TAP_DAC_B = 5'b01110;
    parameter TXPOST_TAP_PD_A = "TRUE";
    parameter TXPOST_TAP_PD_B = "TRUE";
    parameter TXPRE_PRDRV_DAC_A = 3'b111;
    parameter TXPRE_PRDRV_DAC_B = 3'b111;
    parameter TXPRE_TAP_DAC_A = 5'b00000;
    parameter TXPRE_TAP_DAC_B = 5'b00000;
    parameter TXPRE_TAP_PD_A = "TRUE";
    parameter TXPRE_TAP_PD_B = "TRUE";
    parameter TXSLEWRATE_A = "FALSE";
    parameter TXSLEWRATE_B = "FALSE";
    parameter TXTERMTRIM_A = 4'b1100;
    parameter TXTERMTRIM_B = 4'b1100;
    parameter TX_BUFFER_USE_A = "TRUE";
    parameter TX_BUFFER_USE_B = "TRUE";
    parameter TX_CLOCK_DIVIDER_A = 2'b00;
    parameter TX_CLOCK_DIVIDER_B = 2'b00;
    parameter VCODAC_INIT_A = 10'b1010000000;
    parameter VCODAC_INIT_B = 10'b1010000000;
    parameter VCO_CTRL_ENABLE_A = "TRUE";
    parameter VCO_CTRL_ENABLE_B = "TRUE";
    parameter VREFBIASMODE_A = 2'b11;
    parameter VREFBIASMODE_B = 2'b11;
    output DRDYA;
    output DRDYB;
    output RXBUFERRA;
    output RXBUFERRB;
    output RXCALFAILA;
    output RXCALFAILB;
    output RXCOMMADETA;
    output RXCOMMADETB;
    output RXCYCLELIMITA;
    output RXCYCLELIMITB;
    output RXLOCKA;
    output RXLOCKB;
    output RXMCLKA;
    output RXMCLKB;
    output RXPCSHCLKOUTA;
    output RXPCSHCLKOUTB;
    output RXREALIGNA;
    output RXREALIGNB;
    output RXRECCLK1A;
    output RXRECCLK1B;
    output RXRECCLK2A;
    output RXRECCLK2B;
    output RXSIGDETA;
    output RXSIGDETB;
    output TX1NA;
    output TX1NB;
    output TX1PA;
    output TX1PB;
    output TXBUFERRA;
    output TXBUFERRB;
    output TXCALFAILA;
    output TXCALFAILB;
    output TXCYCLELIMITA;
    output TXCYCLELIMITB;
    output TXLOCKA;
    output TXLOCKB;
    output TXOUTCLK1A;
    output TXOUTCLK1B;
    output TXOUTCLK2A;
    output TXOUTCLK2B;
    output TXPCSHCLKOUTA;
    output TXPCSHCLKOUTB;
    output [15:0] DOA;
    output [15:0] DOB;
    output [1:0] RXLOSSOFSYNCA;
    output [1:0] RXLOSSOFSYNCB;
    output [31:0] RXCRCOUTA;
    output [31:0] RXCRCOUTB;
    output [31:0] TXCRCOUTA;
    output [31:0] TXCRCOUTB;
    output [4:0] CHBONDOA;
    output [4:0] CHBONDOB;
    output [5:0] RXSTATUSA;
    output [5:0] RXSTATUSB;
    output [63:0] RXDATAA;
    output [63:0] RXDATAB;
    output [7:0] RXCHARISCOMMAA;
    output [7:0] RXCHARISCOMMAB;
    output [7:0] RXCHARISKA;
    output [7:0] RXCHARISKB;
    output [7:0] RXDISPERRA;
    output [7:0] RXDISPERRB;
    output [7:0] RXNOTINTABLEA;
    output [7:0] RXNOTINTABLEB;
    output [7:0] RXRUNDISPA;
    output [7:0] RXRUNDISPB;
    output [7:0] TXKERRA;
    output [7:0] TXKERRB;
    output [7:0] TXRUNDISPA;
    output [7:0] TXRUNDISPB;
    input DCLKA;
    input DCLKB;
    input DENA;
    input DENB;
    input DWEA;
    input DWEB;
    input ENCHANSYNCA;
    input ENCHANSYNCB;
    input ENMCOMMAALIGNA;
    input ENMCOMMAALIGNB;
    input ENPCOMMAALIGNA;
    input ENPCOMMAALIGNB;
    input GREFCLKA;
    input GREFCLKB;
    input POWERDOWNA;
    input POWERDOWNB;
    input REFCLK1A;
    input REFCLK1B;
    input REFCLK2A;
    input REFCLK2B;
    input RX1NA;
    input RX1NB;
    input RX1PA;
    input RX1PB;
    input RXBLOCKSYNC64B66BUSEA;
    input RXBLOCKSYNC64B66BUSEB;
    input RXCLKSTABLEA;
    input RXCLKSTABLEB;
    input RXCOMMADETUSEA;
    input RXCOMMADETUSEB;
    input RXCRCCLKA;
    input RXCRCCLKB;
    input RXCRCDATAVALIDA;
    input RXCRCDATAVALIDB;
    input RXCRCINITA;
    input RXCRCINITB;
    input RXCRCINTCLKA;
    input RXCRCINTCLKB;
    input RXCRCPDA;
    input RXCRCPDB;
    input RXCRCRESETA;
    input RXCRCRESETB;
    input RXDEC64B66BUSEA;
    input RXDEC64B66BUSEB;
    input RXDEC8B10BUSEA;
    input RXDEC8B10BUSEB;
    input RXDESCRAM64B66BUSEA;
    input RXDESCRAM64B66BUSEB;
    input RXIGNOREBTFA;
    input RXIGNOREBTFB;
    input RXPMARESETA;
    input RXPMARESETB;
    input RXPOLARITYA;
    input RXPOLARITYB;
    input RXRESETA;
    input RXRESETB;
    input RXSLIDEA;
    input RXSLIDEB;
    input RXSYNCA;
    input RXSYNCB;
    input RXUSRCLK2A;
    input RXUSRCLK2B;
    input RXUSRCLKA;
    input RXUSRCLKB;
    input TXCLKSTABLEA;
    input TXCLKSTABLEB;
    input TXCRCCLKA;
    input TXCRCCLKB;
    input TXCRCDATAVALIDA;
    input TXCRCDATAVALIDB;
    input TXCRCINITA;
    input TXCRCINITB;
    input TXCRCINTCLKA;
    input TXCRCINTCLKB;
    input TXCRCPDA;
    input TXCRCPDB;
    input TXCRCRESETA;
    input TXCRCRESETB;
    input TXENC64B66BUSEA;
    input TXENC64B66BUSEB;
    input TXENC8B10BUSEA;
    input TXENC8B10BUSEB;
    input TXENOOBA;
    input TXENOOBB;
    input TXGEARBOX64B66BUSEA;
    input TXGEARBOX64B66BUSEB;
    input TXINHIBITA;
    input TXINHIBITB;
    input TXPMARESETA;
    input TXPMARESETB;
    input TXPOLARITYA;
    input TXPOLARITYB;
    input TXRESETA;
    input TXRESETB;
    input TXSCRAM64B66BUSEA;
    input TXSCRAM64B66BUSEB;
    input TXSYNCA;
    input TXSYNCB;
    input TXUSRCLK2A;
    input TXUSRCLK2B;
    input TXUSRCLKA;
    input TXUSRCLKB;
    input [15:0] DIA;
    input [15:0] DIB;
    input [1:0] LOOPBACKA;
    input [1:0] LOOPBACKB;
    input [1:0] RXDATAWIDTHA;
    input [1:0] RXDATAWIDTHB;
    input [1:0] RXINTDATAWIDTHA;
    input [1:0] RXINTDATAWIDTHB;
    input [1:0] TXDATAWIDTHA;
    input [1:0] TXDATAWIDTHB;
    input [1:0] TXINTDATAWIDTHA;
    input [1:0] TXINTDATAWIDTHB;
    input [2:0] RXCRCDATAWIDTHA;
    input [2:0] RXCRCDATAWIDTHB;
    input [2:0] TXCRCDATAWIDTHA;
    input [2:0] TXCRCDATAWIDTHB;
    input [4:0] CHBONDIA;
    input [4:0] CHBONDIB;
    input [63:0] RXCRCINA;
    input [63:0] RXCRCINB;
    input [63:0] TXCRCINA;
    input [63:0] TXCRCINB;
    input [63:0] TXDATAA;
    input [63:0] TXDATAB;
    input [7:0] DADDRA;
    input [7:0] DADDRB;
    input [7:0] TXBYPASS8B10BA;
    input [7:0] TXBYPASS8B10BB;
    input [7:0] TXCHARDISPMODEA;
    input [7:0] TXCHARDISPMODEB;
    input [7:0] TXCHARDISPVALA;
    input [7:0] TXCHARDISPVALB;
    input [7:0] TXCHARISKA;
    input [7:0] TXCHARISKB;
endmodule

module GT11CLK (...);
    parameter REFCLKSEL = "MGTCLK";
    parameter SYNCLK1OUTEN = "ENABLE";
    parameter SYNCLK2OUTEN = "DISABLE";
    output SYNCLK1OUT;
    output SYNCLK2OUT;
    input MGTCLKN;
    input MGTCLKP;
    input REFCLK;
    input RXBCLK;
    input SYNCLK1IN;
    input SYNCLK2IN;
endmodule

module GT11CLK_MGT (...);
    parameter SYNCLK1OUTEN = "ENABLE";
    parameter SYNCLK2OUTEN = "DISABLE";
    output SYNCLK1OUT;
    output SYNCLK2OUT;
    input MGTCLKN;
    input MGTCLKP;
endmodule

module GTP_DUAL (...);
    parameter AC_CAP_DIS_0 = "TRUE";
    parameter AC_CAP_DIS_1 = "TRUE";
    parameter CHAN_BOND_MODE_0 = "OFF";
    parameter CHAN_BOND_MODE_1 = "OFF";
    parameter CHAN_BOND_SEQ_2_USE_0 = "TRUE";
    parameter CHAN_BOND_SEQ_2_USE_1 = "TRUE";
    parameter CLKINDC_B = "TRUE";
    parameter CLK_CORRECT_USE_0 = "TRUE";
    parameter CLK_CORRECT_USE_1 = "TRUE";
    parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
    parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
    parameter CLK_COR_PRECEDENCE_0 = "TRUE";
    parameter CLK_COR_PRECEDENCE_1 = "TRUE";
    parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
    parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
    parameter COMMA_DOUBLE_0 = "FALSE";
    parameter COMMA_DOUBLE_1 = "FALSE";
    parameter DEC_MCOMMA_DETECT_0 = "TRUE";
    parameter DEC_MCOMMA_DETECT_1 = "TRUE";
    parameter DEC_PCOMMA_DETECT_0 = "TRUE";
    parameter DEC_PCOMMA_DETECT_1 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
    parameter MCOMMA_DETECT_0 = "TRUE";
    parameter MCOMMA_DETECT_1 = "TRUE";
    parameter OVERSAMPLE_MODE = "FALSE";
    parameter PCI_EXPRESS_MODE_0 = "TRUE";
    parameter PCI_EXPRESS_MODE_1 = "TRUE";
    parameter PCOMMA_DETECT_0 = "TRUE";
    parameter PCOMMA_DETECT_1 = "TRUE";
    parameter PLL_SATA_0 = "FALSE";
    parameter PLL_SATA_1 = "FALSE";
    parameter RCV_TERM_GND_0 = "TRUE";
    parameter RCV_TERM_GND_1 = "TRUE";
    parameter RCV_TERM_MID_0 = "FALSE";
    parameter RCV_TERM_MID_1 = "FALSE";
    parameter RCV_TERM_VTTRX_0 = "FALSE";
    parameter RCV_TERM_VTTRX_1 = "FALSE";
    parameter RX_BUFFER_USE_0 = "TRUE";
    parameter RX_BUFFER_USE_1 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
    parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
    parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
    parameter RX_SLIDE_MODE_0 = "PCS";
    parameter RX_SLIDE_MODE_1 = "PCS";
    parameter RX_STATUS_FMT_0 = "PCIE";
    parameter RX_STATUS_FMT_1 = "PCIE";
    parameter RX_XCLK_SEL_0 = "RXREC";
    parameter RX_XCLK_SEL_1 = "RXREC";
    parameter SIM_PLL_PERDIV2 = 9'h190;
    parameter SIM_RECEIVER_DETECT_PASS0 = "FALSE";
    parameter SIM_RECEIVER_DETECT_PASS1 = "FALSE";
    parameter TERMINATION_OVRD = "FALSE";
    parameter TX_BUFFER_USE_0 = "TRUE";
    parameter TX_BUFFER_USE_1 = "TRUE";
    parameter TX_DIFF_BOOST_0 = "TRUE";
    parameter TX_DIFF_BOOST_1 = "TRUE";
    parameter TX_XCLK_SEL_0 = "TXUSR";
    parameter TX_XCLK_SEL_1 = "TXUSR";
    parameter [15:0] TRANS_TIME_FROM_P2_0 = 16'h003c;
    parameter [15:0] TRANS_TIME_FROM_P2_1 = 16'h003c;
    parameter [15:0] TRANS_TIME_NON_P2_0 = 16'h0019;
    parameter [15:0] TRANS_TIME_NON_P2_1 = 16'h0019;
    parameter [15:0] TRANS_TIME_TO_P2_0 = 16'h0064;
    parameter [15:0] TRANS_TIME_TO_P2_1 = 16'h0064;
    parameter [24:0] PMA_RX_CFG_0 = 25'h09f0089;
    parameter [24:0] PMA_RX_CFG_1 = 25'h09f0089;
    parameter [26:0] PMA_CDR_SCAN_0 = 27'h6c07640;
    parameter [26:0] PMA_CDR_SCAN_1 = 27'h6c07640;
    parameter [27:0] PCS_COM_CFG = 28'h1680a0e;
    parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b001;
    parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b001;
    parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
    parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
    parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
    parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
    parameter [31:0] PRBS_ERR_THRESHOLD_0 = 32'h1;
    parameter [31:0] PRBS_ERR_THRESHOLD_1 = 32'h1;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
    parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
    parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
    parameter [4:0] TERMINATION_CTRL = 5'b10100;
    parameter [4:0] TXRX_INVERT_0 = 5'b00000;
    parameter [4:0] TXRX_INVERT_1 = 5'b00000;
    parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
    parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0;
    parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
    parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
    parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
    parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
    parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
    parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
    parameter ALIGN_COMMA_WORD_0 = 1;
    parameter ALIGN_COMMA_WORD_1 = 1;
    parameter CHAN_BOND_1_MAX_SKEW_0 = 7;
    parameter CHAN_BOND_1_MAX_SKEW_1 = 7;
    parameter CHAN_BOND_2_MAX_SKEW_0 = 1;
    parameter CHAN_BOND_2_MAX_SKEW_1 = 1;
    parameter CHAN_BOND_LEVEL_0 = 0;
    parameter CHAN_BOND_LEVEL_1 = 0;
    parameter CHAN_BOND_SEQ_LEN_0 = 4;
    parameter CHAN_BOND_SEQ_LEN_1 = 4;
    parameter CLK25_DIVIDER = 4;
    parameter CLK_COR_ADJ_LEN_0 = 1;
    parameter CLK_COR_ADJ_LEN_1 = 1;
    parameter CLK_COR_DET_LEN_0 = 1;
    parameter CLK_COR_DET_LEN_1 = 1;
    parameter CLK_COR_MAX_LAT_0 = 18;
    parameter CLK_COR_MAX_LAT_1 = 18;
    parameter CLK_COR_MIN_LAT_0 = 16;
    parameter CLK_COR_MIN_LAT_1 = 16;
    parameter CLK_COR_REPEAT_WAIT_0 = 5;
    parameter CLK_COR_REPEAT_WAIT_1 = 5;
    parameter OOB_CLK_DIVIDER = 4;
    parameter PLL_DIVSEL_FB = 5;
    parameter PLL_DIVSEL_REF = 2;
    parameter PLL_RXDIVSEL_OUT_0 = 1;
    parameter PLL_RXDIVSEL_OUT_1 = 1;
    parameter PLL_TXDIVSEL_COMM_OUT = 1;
    parameter PLL_TXDIVSEL_OUT_0 = 1;
    parameter PLL_TXDIVSEL_OUT_1 = 1;
    parameter RX_LOS_INVALID_INCR_0 = 8;
    parameter RX_LOS_INVALID_INCR_1 = 8;
    parameter RX_LOS_THRESHOLD_0 = 128;
    parameter RX_LOS_THRESHOLD_1 = 128;
    parameter SATA_MAX_BURST_0 = 7;
    parameter SATA_MAX_BURST_1 = 7;
    parameter SATA_MAX_INIT_0 = 22;
    parameter SATA_MAX_INIT_1 = 22;
    parameter SATA_MAX_WAKE_0 = 7;
    parameter SATA_MAX_WAKE_1 = 7;
    parameter SATA_MIN_BURST_0 = 4;
    parameter SATA_MIN_BURST_1 = 4;
    parameter SATA_MIN_INIT_0 = 12;
    parameter SATA_MIN_INIT_1 = 12;
    parameter SATA_MIN_WAKE_0 = 4;
    parameter SATA_MIN_WAKE_1 = 4;
    parameter SIM_GTPRESET_SPEEDUP = 0;
    parameter TERMINATION_IMP_0 = 50;
    parameter TERMINATION_IMP_1 = 50;
    parameter TX_SYNC_FILTERB = 1;
    output DRDY;
    output PHYSTATUS0;
    output PHYSTATUS1;
    output PLLLKDET;
    output REFCLKOUT;
    output RESETDONE0;
    output RESETDONE1;
    output RXBYTEISALIGNED0;
    output RXBYTEISALIGNED1;
    output RXBYTEREALIGN0;
    output RXBYTEREALIGN1;
    output RXCHANBONDSEQ0;
    output RXCHANBONDSEQ1;
    output RXCHANISALIGNED0;
    output RXCHANISALIGNED1;
    output RXCHANREALIGN0;
    output RXCHANREALIGN1;
    output RXCOMMADET0;
    output RXCOMMADET1;
    output RXELECIDLE0;
    output RXELECIDLE1;
    output RXOVERSAMPLEERR0;
    output RXOVERSAMPLEERR1;
    output RXPRBSERR0;
    output RXPRBSERR1;
    output RXRECCLK0;
    output RXRECCLK1;
    output RXVALID0;
    output RXVALID1;
    output TXN0;
    output TXN1;
    output TXOUTCLK0;
    output TXOUTCLK1;
    output TXP0;
    output TXP1;
    output [15:0] DO;
    output [15:0] RXDATA0;
    output [15:0] RXDATA1;
    output [1:0] RXCHARISCOMMA0;
    output [1:0] RXCHARISCOMMA1;
    output [1:0] RXCHARISK0;
    output [1:0] RXCHARISK1;
    output [1:0] RXDISPERR0;
    output [1:0] RXDISPERR1;
    output [1:0] RXLOSSOFSYNC0;
    output [1:0] RXLOSSOFSYNC1;
    output [1:0] RXNOTINTABLE0;
    output [1:0] RXNOTINTABLE1;
    output [1:0] RXRUNDISP0;
    output [1:0] RXRUNDISP1;
    output [1:0] TXBUFSTATUS0;
    output [1:0] TXBUFSTATUS1;
    output [1:0] TXKERR0;
    output [1:0] TXKERR1;
    output [1:0] TXRUNDISP0;
    output [1:0] TXRUNDISP1;
    output [2:0] RXBUFSTATUS0;
    output [2:0] RXBUFSTATUS1;
    output [2:0] RXCHBONDO0;
    output [2:0] RXCHBONDO1;
    output [2:0] RXCLKCORCNT0;
    output [2:0] RXCLKCORCNT1;
    output [2:0] RXSTATUS0;
    output [2:0] RXSTATUS1;
    input CLKIN;
    input DCLK;
    input DEN;
    input DWE;
    input GTPRESET;
    input INTDATAWIDTH;
    input PLLLKDETEN;
    input PLLPOWERDOWN;
    input PRBSCNTRESET0;
    input PRBSCNTRESET1;
    input REFCLKPWRDNB;
    input RXBUFRESET0;
    input RXBUFRESET1;
    input RXCDRRESET0;
    input RXCDRRESET1;
    input RXCOMMADETUSE0;
    input RXCOMMADETUSE1;
    input RXDATAWIDTH0;
    input RXDATAWIDTH1;
    input RXDEC8B10BUSE0;
    input RXDEC8B10BUSE1;
    input RXELECIDLERESET0;
    input RXELECIDLERESET1;
    input RXENCHANSYNC0;
    input RXENCHANSYNC1;
    input RXENELECIDLERESETB;
    input RXENEQB0;
    input RXENEQB1;
    input RXENMCOMMAALIGN0;
    input RXENMCOMMAALIGN1;
    input RXENPCOMMAALIGN0;
    input RXENPCOMMAALIGN1;
    input RXENSAMPLEALIGN0;
    input RXENSAMPLEALIGN1;
    input RXN0;
    input RXN1;
    input RXP0;
    input RXP1;
    input RXPMASETPHASE0;
    input RXPMASETPHASE1;
    input RXPOLARITY0;
    input RXPOLARITY1;
    input RXRESET0;
    input RXRESET1;
    input RXSLIDE0;
    input RXSLIDE1;
    input RXUSRCLK0;
    input RXUSRCLK1;
    input RXUSRCLK20;
    input RXUSRCLK21;
    input TXCOMSTART0;
    input TXCOMSTART1;
    input TXCOMTYPE0;
    input TXCOMTYPE1;
    input TXDATAWIDTH0;
    input TXDATAWIDTH1;
    input TXDETECTRX0;
    input TXDETECTRX1;
    input TXELECIDLE0;
    input TXELECIDLE1;
    input TXENC8B10BUSE0;
    input TXENC8B10BUSE1;
    input TXENPMAPHASEALIGN;
    input TXINHIBIT0;
    input TXINHIBIT1;
    input TXPMASETPHASE;
    input TXPOLARITY0;
    input TXPOLARITY1;
    input TXRESET0;
    input TXRESET1;
    input TXUSRCLK0;
    input TXUSRCLK1;
    input TXUSRCLK20;
    input TXUSRCLK21;
    input [15:0] DI;
    input [15:0] TXDATA0;
    input [15:0] TXDATA1;
    input [1:0] RXENPRBSTST0;
    input [1:0] RXENPRBSTST1;
    input [1:0] RXEQMIX0;
    input [1:0] RXEQMIX1;
    input [1:0] RXPOWERDOWN0;
    input [1:0] RXPOWERDOWN1;
    input [1:0] TXBYPASS8B10B0;
    input [1:0] TXBYPASS8B10B1;
    input [1:0] TXCHARDISPMODE0;
    input [1:0] TXCHARDISPMODE1;
    input [1:0] TXCHARDISPVAL0;
    input [1:0] TXCHARDISPVAL1;
    input [1:0] TXCHARISK0;
    input [1:0] TXCHARISK1;
    input [1:0] TXENPRBSTST0;
    input [1:0] TXENPRBSTST1;
    input [1:0] TXPOWERDOWN0;
    input [1:0] TXPOWERDOWN1;
    input [2:0] LOOPBACK0;
    input [2:0] LOOPBACK1;
    input [2:0] RXCHBONDI0;
    input [2:0] RXCHBONDI1;
    input [2:0] TXBUFDIFFCTRL0;
    input [2:0] TXBUFDIFFCTRL1;
    input [2:0] TXDIFFCTRL0;
    input [2:0] TXDIFFCTRL1;
    input [2:0] TXPREEMPHASIS0;
    input [2:0] TXPREEMPHASIS1;
    input [3:0] GTPTEST;
    input [3:0] RXEQPOLE0;
    input [3:0] RXEQPOLE1;
    input [6:0] DADDR;
endmodule

module GTX_DUAL (...);
    parameter STEPPING = "0";
    parameter AC_CAP_DIS_0 = "TRUE";
    parameter AC_CAP_DIS_1 = "TRUE";
    parameter CHAN_BOND_KEEP_ALIGN_0 = "FALSE";
    parameter CHAN_BOND_KEEP_ALIGN_1 = "FALSE";
    parameter CHAN_BOND_MODE_0 = "OFF";
    parameter CHAN_BOND_MODE_1 = "OFF";
    parameter CHAN_BOND_SEQ_2_USE_0 = "TRUE";
    parameter CHAN_BOND_SEQ_2_USE_1 = "TRUE";
    parameter CLKINDC_B = "TRUE";
    parameter CLKRCV_TRST = "FALSE";
    parameter CLK_CORRECT_USE_0 = "TRUE";
    parameter CLK_CORRECT_USE_1 = "TRUE";
    parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
    parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
    parameter CLK_COR_PRECEDENCE_0 = "TRUE";
    parameter CLK_COR_PRECEDENCE_1 = "TRUE";
    parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
    parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
    parameter COMMA_DOUBLE_0 = "FALSE";
    parameter COMMA_DOUBLE_1 = "FALSE";
    parameter DEC_MCOMMA_DETECT_0 = "TRUE";
    parameter DEC_MCOMMA_DETECT_1 = "TRUE";
    parameter DEC_PCOMMA_DETECT_0 = "TRUE";
    parameter DEC_PCOMMA_DETECT_1 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
    parameter MCOMMA_DETECT_0 = "TRUE";
    parameter MCOMMA_DETECT_1 = "TRUE";
    parameter OVERSAMPLE_MODE = "FALSE";
    parameter PCI_EXPRESS_MODE_0 = "TRUE";
    parameter PCI_EXPRESS_MODE_1 = "TRUE";
    parameter PCOMMA_DETECT_0 = "TRUE";
    parameter PCOMMA_DETECT_1 = "TRUE";
    parameter PLL_FB_DCCEN = "FALSE";
    parameter PLL_SATA_0 = "FALSE";
    parameter PLL_SATA_1 = "FALSE";
    parameter RCV_TERM_GND_0 = "TRUE";
    parameter RCV_TERM_GND_1 = "TRUE";
    parameter RCV_TERM_VTTRX_0 = "FALSE";
    parameter RCV_TERM_VTTRX_1 = "FALSE";
    parameter RXGEARBOX_USE_0 = "FALSE";
    parameter RXGEARBOX_USE_1 = "FALSE";
    parameter RX_BUFFER_USE_0 = "TRUE";
    parameter RX_BUFFER_USE_1 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
    parameter RX_EN_IDLE_HOLD_CDR = "FALSE";
    parameter RX_EN_IDLE_HOLD_DFE_0 = "TRUE";
    parameter RX_EN_IDLE_HOLD_DFE_1 = "TRUE";
    parameter RX_EN_IDLE_RESET_BUF_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_BUF_1 = "TRUE";
    parameter RX_EN_IDLE_RESET_FR = "TRUE";
    parameter RX_EN_IDLE_RESET_PH = "TRUE";
    parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
    parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
    parameter RX_SLIDE_MODE_0 = "PCS";
    parameter RX_SLIDE_MODE_1 = "PCS";
    parameter RX_STATUS_FMT_0 = "PCIE";
    parameter RX_STATUS_FMT_1 = "PCIE";
    parameter RX_XCLK_SEL_0 = "RXREC";
    parameter RX_XCLK_SEL_1 = "RXREC";
    parameter SIM_PLL_PERDIV2 = 9'h190;
    parameter SIM_RECEIVER_DETECT_PASS_0 = "FALSE";
    parameter SIM_RECEIVER_DETECT_PASS_1 = "FALSE";
    parameter TERMINATION_OVRD = "FALSE";
    parameter TXGEARBOX_USE_0 = "FALSE";
    parameter TXGEARBOX_USE_1 = "FALSE";
    parameter TX_BUFFER_USE_0 = "TRUE";
    parameter TX_BUFFER_USE_1 = "TRUE";
    parameter TX_XCLK_SEL_0 = "TXUSR";
    parameter TX_XCLK_SEL_1 = "TXUSR";
    parameter [11:0] TRANS_TIME_FROM_P2_0 = 12'h03c;
    parameter [11:0] TRANS_TIME_FROM_P2_1 = 12'h03c;
    parameter [13:0] TX_DETECT_RX_CFG_0 = 14'h1832;
    parameter [13:0] TX_DETECT_RX_CFG_1 = 14'h1832;
    parameter [19:0] PMA_TX_CFG_0 = 20'h00082;
    parameter [19:0] PMA_TX_CFG_1 = 20'h00082;
    parameter [1:0] CM_TRIM_0 = 2'b10;
    parameter [1:0] CM_TRIM_1 = 2'b10;
    parameter [23:0] PLL_COM_CFG = 24'h21680a;
    parameter [24:0] PMA_RX_CFG_0 = 25'h05ce109;
    parameter [24:0] PMA_RX_CFG_1 = 25'h05ce109;
    parameter [26:0] PMA_CDR_SCAN_0 = 27'h6c08040;
    parameter [26:0] PMA_CDR_SCAN_1 = 27'h6c08040;
    parameter [2:0] GEARBOX_ENDEC_0 = 3'b000;
    parameter [2:0] GEARBOX_ENDEC_1 = 3'b000;
    parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b111;
    parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b111;
    parameter [2:0] PLL_LKDET_CFG = 3'b111;
    parameter [2:0] PLL_TDCC_CFG = 3'b000;
    parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
    parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
    parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
    parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
    parameter [2:0] TXRX_INVERT_0 = 3'b000;
    parameter [2:0] TXRX_INVERT_1 = 3'b000;
    parameter [2:0] TX_IDLE_DELAY_0 = 3'b010;
    parameter [2:0] TX_IDLE_DELAY_1 = 3'b010;
    parameter [31:0] PRBS_ERR_THRESHOLD_0 = 32'h1;
    parameter [31:0] PRBS_ERR_THRESHOLD_1 = 32'h1;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
    parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
    parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
    parameter [3:0] RX_IDLE_HI_CNT_0 = 4'b1000;
    parameter [3:0] RX_IDLE_HI_CNT_1 = 4'b1000;
    parameter [3:0] RX_IDLE_LO_CNT_0 = 4'b0000;
    parameter [3:0] RX_IDLE_LO_CNT_1 = 4'b0000;
    parameter [4:0] CDR_PH_ADJ_TIME = 5'b01010;
    parameter [4:0] DFE_CAL_TIME = 5'b00110;
    parameter [4:0] TERMINATION_CTRL = 5'b10100;
    parameter [68:0] PMA_COM_CFG = 69'h0;
    parameter [6:0] PMA_RXSYNC_CFG_0 = 7'h0;
    parameter [6:0] PMA_RXSYNC_CFG_1 = 7'h0;
    parameter [7:0] PLL_CP_CFG = 8'h00;
    parameter [7:0] TRANS_TIME_NON_P2_0 = 8'h19;
    parameter [7:0] TRANS_TIME_NON_P2_1 = 8'h19;
    parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
    parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0;
    parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0;
    parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
    parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
    parameter [9:0] DFE_CFG_0 = 10'b0001111011;
    parameter [9:0] DFE_CFG_1 = 10'b0001111011;
    parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
    parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
    parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
    parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
    parameter [9:0] TRANS_TIME_TO_P2_0 = 10'h064;
    parameter [9:0] TRANS_TIME_TO_P2_1 = 10'h064;
    parameter ALIGN_COMMA_WORD_0 = 1;
    parameter ALIGN_COMMA_WORD_1 = 1;
    parameter CB2_INH_CC_PERIOD_0 = 8;
    parameter CB2_INH_CC_PERIOD_1 = 8;
    parameter CHAN_BOND_1_MAX_SKEW_0 = 7;
    parameter CHAN_BOND_1_MAX_SKEW_1 = 7;
    parameter CHAN_BOND_2_MAX_SKEW_0 = 1;
    parameter CHAN_BOND_2_MAX_SKEW_1 = 1;
    parameter CHAN_BOND_LEVEL_0 = 0;
    parameter CHAN_BOND_LEVEL_1 = 0;
    parameter CHAN_BOND_SEQ_LEN_0 = 4;
    parameter CHAN_BOND_SEQ_LEN_1 = 4;
    parameter CLK25_DIVIDER = 4;
    parameter CLK_COR_ADJ_LEN_0 = 1;
    parameter CLK_COR_ADJ_LEN_1 = 1;
    parameter CLK_COR_DET_LEN_0 = 1;
    parameter CLK_COR_DET_LEN_1 = 1;
    parameter CLK_COR_MAX_LAT_0 = 18;
    parameter CLK_COR_MAX_LAT_1 = 18;
    parameter CLK_COR_MIN_LAT_0 = 16;
    parameter CLK_COR_MIN_LAT_1 = 16;
    parameter CLK_COR_REPEAT_WAIT_0 = 5;
    parameter CLK_COR_REPEAT_WAIT_1 = 5;
    parameter OOB_CLK_DIVIDER = 4;
    parameter PLL_DIVSEL_FB = 5;
    parameter PLL_DIVSEL_REF = 2;
    parameter PLL_RXDIVSEL_OUT_0 = 1;
    parameter PLL_RXDIVSEL_OUT_1 = 1;
    parameter PLL_TXDIVSEL_OUT_0 = 1;
    parameter PLL_TXDIVSEL_OUT_1 = 1;
    parameter RX_LOS_INVALID_INCR_0 = 8;
    parameter RX_LOS_INVALID_INCR_1 = 8;
    parameter RX_LOS_THRESHOLD_0 = 128;
    parameter RX_LOS_THRESHOLD_1 = 128;
    parameter SATA_MAX_BURST_0 = 7;
    parameter SATA_MAX_BURST_1 = 7;
    parameter SATA_MAX_INIT_0 = 22;
    parameter SATA_MAX_INIT_1 = 22;
    parameter SATA_MAX_WAKE_0 = 7;
    parameter SATA_MAX_WAKE_1 = 7;
    parameter SATA_MIN_BURST_0 = 4;
    parameter SATA_MIN_BURST_1 = 4;
    parameter SATA_MIN_INIT_0 = 12;
    parameter SATA_MIN_INIT_1 = 12;
    parameter SATA_MIN_WAKE_0 = 4;
    parameter SATA_MIN_WAKE_1 = 4;
    parameter SIM_GTXRESET_SPEEDUP = 0;
    parameter TERMINATION_IMP_0 = 50;
    parameter TERMINATION_IMP_1 = 50;
    output DRDY;
    output PHYSTATUS0;
    output PHYSTATUS1;
    output PLLLKDET;
    output REFCLKOUT;
    output RESETDONE0;
    output RESETDONE1;
    output RXBYTEISALIGNED0;
    output RXBYTEISALIGNED1;
    output RXBYTEREALIGN0;
    output RXBYTEREALIGN1;
    output RXCHANBONDSEQ0;
    output RXCHANBONDSEQ1;
    output RXCHANISALIGNED0;
    output RXCHANISALIGNED1;
    output RXCHANREALIGN0;
    output RXCHANREALIGN1;
    output RXCOMMADET0;
    output RXCOMMADET1;
    output RXDATAVALID0;
    output RXDATAVALID1;
    output RXELECIDLE0;
    output RXELECIDLE1;
    output RXHEADERVALID0;
    output RXHEADERVALID1;
    output RXOVERSAMPLEERR0;
    output RXOVERSAMPLEERR1;
    output RXPRBSERR0;
    output RXPRBSERR1;
    output RXRECCLK0;
    output RXRECCLK1;
    output RXSTARTOFSEQ0;
    output RXSTARTOFSEQ1;
    output RXVALID0;
    output RXVALID1;
    output TXGEARBOXREADY0;
    output TXGEARBOXREADY1;
    output TXN0;
    output TXN1;
    output TXOUTCLK0;
    output TXOUTCLK1;
    output TXP0;
    output TXP1;
    output [15:0] DO;
    output [1:0] RXLOSSOFSYNC0;
    output [1:0] RXLOSSOFSYNC1;
    output [1:0] TXBUFSTATUS0;
    output [1:0] TXBUFSTATUS1;
    output [2:0] DFESENSCAL0;
    output [2:0] DFESENSCAL1;
    output [2:0] RXBUFSTATUS0;
    output [2:0] RXBUFSTATUS1;
    output [2:0] RXCLKCORCNT0;
    output [2:0] RXCLKCORCNT1;
    output [2:0] RXHEADER0;
    output [2:0] RXHEADER1;
    output [2:0] RXSTATUS0;
    output [2:0] RXSTATUS1;
    output [31:0] RXDATA0;
    output [31:0] RXDATA1;
    output [3:0] DFETAP3MONITOR0;
    output [3:0] DFETAP3MONITOR1;
    output [3:0] DFETAP4MONITOR0;
    output [3:0] DFETAP4MONITOR1;
    output [3:0] RXCHARISCOMMA0;
    output [3:0] RXCHARISCOMMA1;
    output [3:0] RXCHARISK0;
    output [3:0] RXCHARISK1;
    output [3:0] RXCHBONDO0;
    output [3:0] RXCHBONDO1;
    output [3:0] RXDISPERR0;
    output [3:0] RXDISPERR1;
    output [3:0] RXNOTINTABLE0;
    output [3:0] RXNOTINTABLE1;
    output [3:0] RXRUNDISP0;
    output [3:0] RXRUNDISP1;
    output [3:0] TXKERR0;
    output [3:0] TXKERR1;
    output [3:0] TXRUNDISP0;
    output [3:0] TXRUNDISP1;
    output [4:0] DFEEYEDACMONITOR0;
    output [4:0] DFEEYEDACMONITOR1;
    output [4:0] DFETAP1MONITOR0;
    output [4:0] DFETAP1MONITOR1;
    output [4:0] DFETAP2MONITOR0;
    output [4:0] DFETAP2MONITOR1;
    output [5:0] DFECLKDLYADJMONITOR0;
    output [5:0] DFECLKDLYADJMONITOR1;
    input CLKIN;
    input DCLK;
    input DEN;
    input DWE;
    input GTXRESET;
    input INTDATAWIDTH;
    input PLLLKDETEN;
    input PLLPOWERDOWN;
    input PRBSCNTRESET0;
    input PRBSCNTRESET1;
    input REFCLKPWRDNB;
    input RXBUFRESET0;
    input RXBUFRESET1;
    input RXCDRRESET0;
    input RXCDRRESET1;
    input RXCOMMADETUSE0;
    input RXCOMMADETUSE1;
    input RXDEC8B10BUSE0;
    input RXDEC8B10BUSE1;
    input RXENCHANSYNC0;
    input RXENCHANSYNC1;
    input RXENEQB0;
    input RXENEQB1;
    input RXENMCOMMAALIGN0;
    input RXENMCOMMAALIGN1;
    input RXENPCOMMAALIGN0;
    input RXENPCOMMAALIGN1;
    input RXENPMAPHASEALIGN0;
    input RXENPMAPHASEALIGN1;
    input RXENSAMPLEALIGN0;
    input RXENSAMPLEALIGN1;
    input RXGEARBOXSLIP0;
    input RXGEARBOXSLIP1;
    input RXN0;
    input RXN1;
    input RXP0;
    input RXP1;
    input RXPMASETPHASE0;
    input RXPMASETPHASE1;
    input RXPOLARITY0;
    input RXPOLARITY1;
    input RXRESET0;
    input RXRESET1;
    input RXSLIDE0;
    input RXSLIDE1;
    input RXUSRCLK0;
    input RXUSRCLK1;
    input RXUSRCLK20;
    input RXUSRCLK21;
    input TXCOMSTART0;
    input TXCOMSTART1;
    input TXCOMTYPE0;
    input TXCOMTYPE1;
    input TXDETECTRX0;
    input TXDETECTRX1;
    input TXELECIDLE0;
    input TXELECIDLE1;
    input TXENC8B10BUSE0;
    input TXENC8B10BUSE1;
    input TXENPMAPHASEALIGN0;
    input TXENPMAPHASEALIGN1;
    input TXINHIBIT0;
    input TXINHIBIT1;
    input TXPMASETPHASE0;
    input TXPMASETPHASE1;
    input TXPOLARITY0;
    input TXPOLARITY1;
    input TXRESET0;
    input TXRESET1;
    input TXSTARTSEQ0;
    input TXSTARTSEQ1;
    input TXUSRCLK0;
    input TXUSRCLK1;
    input TXUSRCLK20;
    input TXUSRCLK21;
    input [13:0] GTXTEST;
    input [15:0] DI;
    input [1:0] RXDATAWIDTH0;
    input [1:0] RXDATAWIDTH1;
    input [1:0] RXENPRBSTST0;
    input [1:0] RXENPRBSTST1;
    input [1:0] RXEQMIX0;
    input [1:0] RXEQMIX1;
    input [1:0] RXPOWERDOWN0;
    input [1:0] RXPOWERDOWN1;
    input [1:0] TXDATAWIDTH0;
    input [1:0] TXDATAWIDTH1;
    input [1:0] TXENPRBSTST0;
    input [1:0] TXENPRBSTST1;
    input [1:0] TXPOWERDOWN0;
    input [1:0] TXPOWERDOWN1;
    input [2:0] LOOPBACK0;
    input [2:0] LOOPBACK1;
    input [2:0] TXBUFDIFFCTRL0;
    input [2:0] TXBUFDIFFCTRL1;
    input [2:0] TXDIFFCTRL0;
    input [2:0] TXDIFFCTRL1;
    input [2:0] TXHEADER0;
    input [2:0] TXHEADER1;
    input [31:0] TXDATA0;
    input [31:0] TXDATA1;
    input [3:0] DFETAP30;
    input [3:0] DFETAP31;
    input [3:0] DFETAP40;
    input [3:0] DFETAP41;
    input [3:0] RXCHBONDI0;
    input [3:0] RXCHBONDI1;
    input [3:0] RXEQPOLE0;
    input [3:0] RXEQPOLE1;
    input [3:0] TXBYPASS8B10B0;
    input [3:0] TXBYPASS8B10B1;
    input [3:0] TXCHARDISPMODE0;
    input [3:0] TXCHARDISPMODE1;
    input [3:0] TXCHARDISPVAL0;
    input [3:0] TXCHARDISPVAL1;
    input [3:0] TXCHARISK0;
    input [3:0] TXCHARISK1;
    input [3:0] TXPREEMPHASIS0;
    input [3:0] TXPREEMPHASIS1;
    input [4:0] DFETAP10;
    input [4:0] DFETAP11;
    input [4:0] DFETAP20;
    input [4:0] DFETAP21;
    input [5:0] DFECLKDLYADJ0;
    input [5:0] DFECLKDLYADJ1;
    input [6:0] DADDR;
    input [6:0] TXSEQUENCE0;
    input [6:0] TXSEQUENCE1;
endmodule

module CRC32 (...);
    parameter CRC_INIT = 32'hFFFFFFFF;
    output [31:0] CRCOUT;
    (* clkbuf_sink *)
    input CRCCLK;
    input CRCDATAVALID;
    input [2:0] CRCDATAWIDTH;
    input [31:0] CRCIN;
    input CRCRESET;
endmodule

module CRC64 (...);
    parameter CRC_INIT = 32'hFFFFFFFF;
    output [31:0] CRCOUT;
    (* clkbuf_sink *)
    input CRCCLK;
    input CRCDATAVALID;
    input [2:0] CRCDATAWIDTH;
    input [63:0] CRCIN;
    input CRCRESET;
endmodule

module GTHE1_QUAD (...);
    parameter [15:0] BER_CONST_PTRN0 = 16'h0000;
    parameter [15:0] BER_CONST_PTRN1 = 16'h0000;
    parameter [15:0] BUFFER_CONFIG_LANE0 = 16'h4004;
    parameter [15:0] BUFFER_CONFIG_LANE1 = 16'h4004;
    parameter [15:0] BUFFER_CONFIG_LANE2 = 16'h4004;
    parameter [15:0] BUFFER_CONFIG_LANE3 = 16'h4004;
    parameter [15:0] DFE_TRAIN_CTRL_LANE0 = 16'h0000;
    parameter [15:0] DFE_TRAIN_CTRL_LANE1 = 16'h0000;
    parameter [15:0] DFE_TRAIN_CTRL_LANE2 = 16'h0000;
    parameter [15:0] DFE_TRAIN_CTRL_LANE3 = 16'h0000;
    parameter [15:0] DLL_CFG0 = 16'h8202;
    parameter [15:0] DLL_CFG1 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE3 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE3 = 16'h0000;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE0 = 16'h0002;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE1 = 16'h0002;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE2 = 16'h0002;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE3 = 16'h0002;
    parameter [15:0] E10GBASEKX_CTRL_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEKX_CTRL_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEKX_CTRL_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEKX_CTRL_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_CFG_LANE0 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_CFG_LANE1 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_CFG_LANE2 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_CFG_LANE3 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE0 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE1 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE2 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE3 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE0 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE1 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE2 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE3 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE3 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE3 = 16'h0000;
    parameter [15:0] GLBL0_NOISE_CTRL = 16'hF0B8;
    parameter [15:0] GLBL_AMON_SEL = 16'h0000;
    parameter [15:0] GLBL_DMON_SEL = 16'h0200;
    parameter [15:0] GLBL_PWR_CTRL = 16'h0000;
    parameter [0:0] GTH_CFG_PWRUP_LANE0 = 1'b1;
    parameter [0:0] GTH_CFG_PWRUP_LANE1 = 1'b1;
    parameter [0:0] GTH_CFG_PWRUP_LANE2 = 1'b1;
    parameter [0:0] GTH_CFG_PWRUP_LANE3 = 1'b1;
    parameter [15:0] LANE_AMON_SEL = 16'h00F0;
    parameter [15:0] LANE_DMON_SEL = 16'h0000;
    parameter [15:0] LANE_LNK_CFGOVRD = 16'h0000;
    parameter [15:0] LANE_PWR_CTRL_LANE0 = 16'h0400;
    parameter [15:0] LANE_PWR_CTRL_LANE1 = 16'h0400;
    parameter [15:0] LANE_PWR_CTRL_LANE2 = 16'h0400;
    parameter [15:0] LANE_PWR_CTRL_LANE3 = 16'h0400;
    parameter [15:0] LNK_TRN_CFG_LANE0 = 16'h0000;
    parameter [15:0] LNK_TRN_CFG_LANE1 = 16'h0000;
    parameter [15:0] LNK_TRN_CFG_LANE2 = 16'h0000;
    parameter [15:0] LNK_TRN_CFG_LANE3 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE0 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE1 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE2 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE3 = 16'h0000;
    parameter [15:0] MISC_CFG = 16'h0008;
    parameter [15:0] MODE_CFG1 = 16'h0000;
    parameter [15:0] MODE_CFG2 = 16'h0000;
    parameter [15:0] MODE_CFG3 = 16'h0000;
    parameter [15:0] MODE_CFG4 = 16'h0000;
    parameter [15:0] MODE_CFG5 = 16'h0000;
    parameter [15:0] MODE_CFG6 = 16'h0000;
    parameter [15:0] MODE_CFG7 = 16'h0000;
    parameter [15:0] PCS_ABILITY_LANE0 = 16'h0010;
    parameter [15:0] PCS_ABILITY_LANE1 = 16'h0010;
    parameter [15:0] PCS_ABILITY_LANE2 = 16'h0010;
    parameter [15:0] PCS_ABILITY_LANE3 = 16'h0010;
    parameter [15:0] PCS_CTRL1_LANE0 = 16'h2040;
    parameter [15:0] PCS_CTRL1_LANE1 = 16'h2040;
    parameter [15:0] PCS_CTRL1_LANE2 = 16'h2040;
    parameter [15:0] PCS_CTRL1_LANE3 = 16'h2040;
    parameter [15:0] PCS_CTRL2_LANE0 = 16'h0000;
    parameter [15:0] PCS_CTRL2_LANE1 = 16'h0000;
    parameter [15:0] PCS_CTRL2_LANE2 = 16'h0000;
    parameter [15:0] PCS_CTRL2_LANE3 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_0_LANE0 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_0_LANE1 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_0_LANE2 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_0_LANE3 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_1_LANE0 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_1_LANE1 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_1_LANE2 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_1_LANE3 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE0 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE1 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE2 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE3 = 16'h0000;
    parameter [15:0] PCS_RESET_1_LANE0 = 16'h0002;
    parameter [15:0] PCS_RESET_1_LANE1 = 16'h0002;
    parameter [15:0] PCS_RESET_1_LANE2 = 16'h0002;
    parameter [15:0] PCS_RESET_1_LANE3 = 16'h0002;
    parameter [15:0] PCS_RESET_LANE0 = 16'h0000;
    parameter [15:0] PCS_RESET_LANE1 = 16'h0000;
    parameter [15:0] PCS_RESET_LANE2 = 16'h0000;
    parameter [15:0] PCS_RESET_LANE3 = 16'h0000;
    parameter [15:0] PCS_TYPE_LANE0 = 16'h002C;
    parameter [15:0] PCS_TYPE_LANE1 = 16'h002C;
    parameter [15:0] PCS_TYPE_LANE2 = 16'h002C;
    parameter [15:0] PCS_TYPE_LANE3 = 16'h002C;
    parameter [15:0] PLL_CFG0 = 16'h95DF;
    parameter [15:0] PLL_CFG1 = 16'h81C0;
    parameter [15:0] PLL_CFG2 = 16'h0424;
    parameter [15:0] PMA_CTRL1_LANE0 = 16'h0000;
    parameter [15:0] PMA_CTRL1_LANE1 = 16'h0000;
    parameter [15:0] PMA_CTRL1_LANE2 = 16'h0000;
    parameter [15:0] PMA_CTRL1_LANE3 = 16'h0000;
    parameter [15:0] PMA_CTRL2_LANE0 = 16'h000B;
    parameter [15:0] PMA_CTRL2_LANE1 = 16'h000B;
    parameter [15:0] PMA_CTRL2_LANE2 = 16'h000B;
    parameter [15:0] PMA_CTRL2_LANE3 = 16'h000B;
    parameter [15:0] PMA_LPBK_CTRL_LANE0 = 16'h0004;
    parameter [15:0] PMA_LPBK_CTRL_LANE1 = 16'h0004;
    parameter [15:0] PMA_LPBK_CTRL_LANE2 = 16'h0004;
    parameter [15:0] PMA_LPBK_CTRL_LANE3 = 16'h0004;
    parameter [15:0] PRBS_BER_CFG0_LANE0 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG0_LANE1 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG0_LANE2 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG0_LANE3 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE0 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE1 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE2 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE3 = 16'h0000;
    parameter [15:0] PRBS_CFG_LANE0 = 16'h000A;
    parameter [15:0] PRBS_CFG_LANE1 = 16'h000A;
    parameter [15:0] PRBS_CFG_LANE2 = 16'h000A;
    parameter [15:0] PRBS_CFG_LANE3 = 16'h000A;
    parameter [15:0] PTRN_CFG0_LSB = 16'h5555;
    parameter [15:0] PTRN_CFG0_MSB = 16'h5555;
    parameter [15:0] PTRN_LEN_CFG = 16'h001F;
    parameter [15:0] PWRUP_DLY = 16'h0000;
    parameter [15:0] RX_AEQ_VAL0_LANE0 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL0_LANE1 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL0_LANE2 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL0_LANE3 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL1_LANE0 = 16'h0000;
    parameter [15:0] RX_AEQ_VAL1_LANE1 = 16'h0000;
    parameter [15:0] RX_AEQ_VAL1_LANE2 = 16'h0000;
    parameter [15:0] RX_AEQ_VAL1_LANE3 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE0 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE1 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE2 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE3 = 16'h0000;
    parameter [15:0] RX_CDR_CTRL0_LANE0 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL0_LANE1 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL0_LANE2 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL0_LANE3 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL1_LANE0 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL1_LANE1 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL1_LANE2 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL1_LANE3 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL2_LANE0 = 16'h2000;
    parameter [15:0] RX_CDR_CTRL2_LANE1 = 16'h2000;
    parameter [15:0] RX_CDR_CTRL2_LANE2 = 16'h2000;
    parameter [15:0] RX_CDR_CTRL2_LANE3 = 16'h2000;
    parameter [15:0] RX_CFG0_LANE0 = 16'h0500;
    parameter [15:0] RX_CFG0_LANE1 = 16'h0500;
    parameter [15:0] RX_CFG0_LANE2 = 16'h0500;
    parameter [15:0] RX_CFG0_LANE3 = 16'h0500;
    parameter [15:0] RX_CFG1_LANE0 = 16'h821F;
    parameter [15:0] RX_CFG1_LANE1 = 16'h821F;
    parameter [15:0] RX_CFG1_LANE2 = 16'h821F;
    parameter [15:0] RX_CFG1_LANE3 = 16'h821F;
    parameter [15:0] RX_CFG2_LANE0 = 16'h1001;
    parameter [15:0] RX_CFG2_LANE1 = 16'h1001;
    parameter [15:0] RX_CFG2_LANE2 = 16'h1001;
    parameter [15:0] RX_CFG2_LANE3 = 16'h1001;
    parameter [15:0] RX_CTLE_CTRL_LANE0 = 16'h008F;
    parameter [15:0] RX_CTLE_CTRL_LANE1 = 16'h008F;
    parameter [15:0] RX_CTLE_CTRL_LANE2 = 16'h008F;
    parameter [15:0] RX_CTLE_CTRL_LANE3 = 16'h008F;
    parameter [15:0] RX_CTRL_OVRD_LANE0 = 16'h000C;
    parameter [15:0] RX_CTRL_OVRD_LANE1 = 16'h000C;
    parameter [15:0] RX_CTRL_OVRD_LANE2 = 16'h000C;
    parameter [15:0] RX_CTRL_OVRD_LANE3 = 16'h000C;
    parameter integer RX_FABRIC_WIDTH0 = 6466;
    parameter integer RX_FABRIC_WIDTH1 = 6466;
    parameter integer RX_FABRIC_WIDTH2 = 6466;
    parameter integer RX_FABRIC_WIDTH3 = 6466;
    parameter [15:0] RX_LOOP_CTRL_LANE0 = 16'h007F;
    parameter [15:0] RX_LOOP_CTRL_LANE1 = 16'h007F;
    parameter [15:0] RX_LOOP_CTRL_LANE2 = 16'h007F;
    parameter [15:0] RX_LOOP_CTRL_LANE3 = 16'h007F;
    parameter [15:0] RX_MVAL0_LANE0 = 16'h0000;
    parameter [15:0] RX_MVAL0_LANE1 = 16'h0000;
    parameter [15:0] RX_MVAL0_LANE2 = 16'h0000;
    parameter [15:0] RX_MVAL0_LANE3 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE0 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE1 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE2 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE3 = 16'h0000;
    parameter [15:0] RX_P0S_CTRL = 16'h1206;
    parameter [15:0] RX_P0_CTRL = 16'h11F0;
    parameter [15:0] RX_P1_CTRL = 16'h120F;
    parameter [15:0] RX_P2_CTRL = 16'h0E0F;
    parameter [15:0] RX_PI_CTRL0 = 16'hD2F0;
    parameter [15:0] RX_PI_CTRL1 = 16'h0080;
    parameter integer SIM_GTHRESET_SPEEDUP = 1;
    parameter SIM_VERSION = "1.0";
    parameter [15:0] SLICE_CFG = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_0_LANE01 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_0_LANE23 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_1_LANE01 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_1_LANE23 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_2_LANE01 = 16'h7FFF;
    parameter [15:0] SLICE_NOISE_CTRL_2_LANE23 = 16'h7FFF;
    parameter [15:0] SLICE_TX_RESET_LANE01 = 16'h0000;
    parameter [15:0] SLICE_TX_RESET_LANE23 = 16'h0000;
    parameter [15:0] TERM_CTRL_LANE0 = 16'h5007;
    parameter [15:0] TERM_CTRL_LANE1 = 16'h5007;
    parameter [15:0] TERM_CTRL_LANE2 = 16'h5007;
    parameter [15:0] TERM_CTRL_LANE3 = 16'h5007;
    parameter [15:0] TX_CFG0_LANE0 = 16'h203D;
    parameter [15:0] TX_CFG0_LANE1 = 16'h203D;
    parameter [15:0] TX_CFG0_LANE2 = 16'h203D;
    parameter [15:0] TX_CFG0_LANE3 = 16'h203D;
    parameter [15:0] TX_CFG1_LANE0 = 16'h0F00;
    parameter [15:0] TX_CFG1_LANE1 = 16'h0F00;
    parameter [15:0] TX_CFG1_LANE2 = 16'h0F00;
    parameter [15:0] TX_CFG1_LANE3 = 16'h0F00;
    parameter [15:0] TX_CFG2_LANE0 = 16'h0081;
    parameter [15:0] TX_CFG2_LANE1 = 16'h0081;
    parameter [15:0] TX_CFG2_LANE2 = 16'h0081;
    parameter [15:0] TX_CFG2_LANE3 = 16'h0081;
    parameter [15:0] TX_CLK_SEL0_LANE0 = 16'h2121;
    parameter [15:0] TX_CLK_SEL0_LANE1 = 16'h2121;
    parameter [15:0] TX_CLK_SEL0_LANE2 = 16'h2121;
    parameter [15:0] TX_CLK_SEL0_LANE3 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE0 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE1 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE2 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE3 = 16'h2121;
    parameter [15:0] TX_DISABLE_LANE0 = 16'h0000;
    parameter [15:0] TX_DISABLE_LANE1 = 16'h0000;
    parameter [15:0] TX_DISABLE_LANE2 = 16'h0000;
    parameter [15:0] TX_DISABLE_LANE3 = 16'h0000;
    parameter integer TX_FABRIC_WIDTH0 = 6466;
    parameter integer TX_FABRIC_WIDTH1 = 6466;
    parameter integer TX_FABRIC_WIDTH2 = 6466;
    parameter integer TX_FABRIC_WIDTH3 = 6466;
    parameter [15:0] TX_P0P0S_CTRL = 16'h060C;
    parameter [15:0] TX_P1P2_CTRL = 16'h0C39;
    parameter [15:0] TX_PREEMPH_LANE0 = 16'h00A1;
    parameter [15:0] TX_PREEMPH_LANE1 = 16'h00A1;
    parameter [15:0] TX_PREEMPH_LANE2 = 16'h00A1;
    parameter [15:0] TX_PREEMPH_LANE3 = 16'h00A1;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE0 = 16'h0060;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE1 = 16'h0060;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE2 = 16'h0060;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE3 = 16'h0060;
    output DRDY;
    output GTHINITDONE;
    output MGMTPCSRDACK;
    output RXCTRLACK0;
    output RXCTRLACK1;
    output RXCTRLACK2;
    output RXCTRLACK3;
    output RXDATATAP0;
    output RXDATATAP1;
    output RXDATATAP2;
    output RXDATATAP3;
    output RXPCSCLKSMPL0;
    output RXPCSCLKSMPL1;
    output RXPCSCLKSMPL2;
    output RXPCSCLKSMPL3;
    output RXUSERCLKOUT0;
    output RXUSERCLKOUT1;
    output RXUSERCLKOUT2;
    output RXUSERCLKOUT3;
    output TSTPATH;
    output TSTREFCLKFAB;
    output TSTREFCLKOUT;
    output TXCTRLACK0;
    output TXCTRLACK1;
    output TXCTRLACK2;
    output TXCTRLACK3;
    output TXDATATAP10;
    output TXDATATAP11;
    output TXDATATAP12;
    output TXDATATAP13;
    output TXDATATAP20;
    output TXDATATAP21;
    output TXDATATAP22;
    output TXDATATAP23;
    output TXN0;
    output TXN1;
    output TXN2;
    output TXN3;
    output TXP0;
    output TXP1;
    output TXP2;
    output TXP3;
    output TXPCSCLKSMPL0;
    output TXPCSCLKSMPL1;
    output TXPCSCLKSMPL2;
    output TXPCSCLKSMPL3;
    output TXUSERCLKOUT0;
    output TXUSERCLKOUT1;
    output TXUSERCLKOUT2;
    output TXUSERCLKOUT3;
    output [15:0] DRPDO;
    output [15:0] MGMTPCSRDDATA;
    output [63:0] RXDATA0;
    output [63:0] RXDATA1;
    output [63:0] RXDATA2;
    output [63:0] RXDATA3;
    output [7:0] RXCODEERR0;
    output [7:0] RXCODEERR1;
    output [7:0] RXCODEERR2;
    output [7:0] RXCODEERR3;
    output [7:0] RXCTRL0;
    output [7:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [7:0] RXDISPERR0;
    output [7:0] RXDISPERR1;
    output [7:0] RXDISPERR2;
    output [7:0] RXDISPERR3;
    output [7:0] RXVALID0;
    output [7:0] RXVALID1;
    output [7:0] RXVALID2;
    output [7:0] RXVALID3;
    input DCLK;
    input DEN;
    input DFETRAINCTRL0;
    input DFETRAINCTRL1;
    input DFETRAINCTRL2;
    input DFETRAINCTRL3;
    input DISABLEDRP;
    input DWE;
    input GTHINIT;
    input GTHRESET;
    input GTHX2LANE01;
    input GTHX2LANE23;
    input GTHX4LANE;
    input MGMTPCSREGRD;
    input MGMTPCSREGWR;
    input POWERDOWN0;
    input POWERDOWN1;
    input POWERDOWN2;
    input POWERDOWN3;
    input REFCLK;
    input RXBUFRESET0;
    input RXBUFRESET1;
    input RXBUFRESET2;
    input RXBUFRESET3;
    input RXENCOMMADET0;
    input RXENCOMMADET1;
    input RXENCOMMADET2;
    input RXENCOMMADET3;
    input RXN0;
    input RXN1;
    input RXN2;
    input RXN3;
    input RXP0;
    input RXP1;
    input RXP2;
    input RXP3;
    input RXPOLARITY0;
    input RXPOLARITY1;
    input RXPOLARITY2;
    input RXPOLARITY3;
    input RXSLIP0;
    input RXSLIP1;
    input RXSLIP2;
    input RXSLIP3;
    input RXUSERCLKIN0;
    input RXUSERCLKIN1;
    input RXUSERCLKIN2;
    input RXUSERCLKIN3;
    input TXBUFRESET0;
    input TXBUFRESET1;
    input TXBUFRESET2;
    input TXBUFRESET3;
    input TXDEEMPH0;
    input TXDEEMPH1;
    input TXDEEMPH2;
    input TXDEEMPH3;
    input TXUSERCLKIN0;
    input TXUSERCLKIN1;
    input TXUSERCLKIN2;
    input TXUSERCLKIN3;
    input [15:0] DADDR;
    input [15:0] DI;
    input [15:0] MGMTPCSREGADDR;
    input [15:0] MGMTPCSWRDATA;
    input [1:0] RXPOWERDOWN0;
    input [1:0] RXPOWERDOWN1;
    input [1:0] RXPOWERDOWN2;
    input [1:0] RXPOWERDOWN3;
    input [1:0] RXRATE0;
    input [1:0] RXRATE1;
    input [1:0] RXRATE2;
    input [1:0] RXRATE3;
    input [1:0] TXPOWERDOWN0;
    input [1:0] TXPOWERDOWN1;
    input [1:0] TXPOWERDOWN2;
    input [1:0] TXPOWERDOWN3;
    input [1:0] TXRATE0;
    input [1:0] TXRATE1;
    input [1:0] TXRATE2;
    input [1:0] TXRATE3;
    input [2:0] PLLREFCLKSEL;
    input [2:0] SAMPLERATE0;
    input [2:0] SAMPLERATE1;
    input [2:0] SAMPLERATE2;
    input [2:0] SAMPLERATE3;
    input [2:0] TXMARGIN0;
    input [2:0] TXMARGIN1;
    input [2:0] TXMARGIN2;
    input [2:0] TXMARGIN3;
    input [3:0] MGMTPCSLANESEL;
    input [4:0] MGMTPCSMMDADDR;
    input [5:0] PLLPCSCLKDIV;
    input [63:0] TXDATA0;
    input [63:0] TXDATA1;
    input [63:0] TXDATA2;
    input [63:0] TXDATA3;
    input [7:0] TXCTRL0;
    input [7:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [7:0] TXCTRL3;
    input [7:0] TXDATAMSB0;
    input [7:0] TXDATAMSB1;
    input [7:0] TXDATAMSB2;
    input [7:0] TXDATAMSB3;
endmodule

module GTXE1 (...);
    parameter AC_CAP_DIS = "TRUE";
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter [1:0] BGTEST_CFG = 2'b00;
    parameter [16:0] BIAS_CFG = 17'h00000;
    parameter [4:0] CDR_PH_ADJ_TIME = 5'b10100;
    parameter integer CHAN_BOND_1_MAX_SKEW = 7;
    parameter integer CHAN_BOND_2_MAX_SKEW = 1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0110111100;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100111100;
    parameter [4:0] CHAN_BOND_SEQ_2_CFG = 5'b00000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter integer CLK_COR_ADJ_LEN = 1;
    parameter integer CLK_COR_DET_LEN = 1;
    parameter CLK_COR_INSERT_IDLE_FLAG = "FALSE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter [1:0] CM_TRIM = 2'b01;
    parameter [9:0] COMMA_10B_ENABLE = 10'b1111111111;
    parameter COMMA_DOUBLE = "FALSE";
    parameter [3:0] COM_BURST_VAL = 4'b1111;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [4:0] DFE_CAL_TIME = 5'b01100;
    parameter [7:0] DFE_CFG = 8'b00011011;
    parameter [2:0] GEARBOX_ENDEC = 3'b000;
    parameter GEN_RXUSRCLK = "TRUE";
    parameter GEN_TXUSRCLK = "TRUE";
    parameter GTX_CFG_PWRUP = "TRUE";
    parameter [9:0] MCOMMA_10B_VALUE = 10'b1010000011;
    parameter MCOMMA_DETECT = "TRUE";
    parameter [2:0] OOBDETECT_THRESHOLD = 3'b011;
    parameter PCI_EXPRESS_MODE = "FALSE";
    parameter [9:0] PCOMMA_10B_VALUE = 10'b0101111100;
    parameter PCOMMA_DETECT = "TRUE";
    parameter PMA_CAS_CLK_EN = "FALSE";
    parameter [26:0] PMA_CDR_SCAN = 27'h640404C;
    parameter [75:0] PMA_CFG = 76'h0040000040000000003;
    parameter [6:0] PMA_RXSYNC_CFG = 7'h00;
    parameter [24:0] PMA_RX_CFG = 25'h05CE048;
    parameter [19:0] PMA_TX_CFG = 20'h00082;
    parameter [9:0] POWER_SAVE = 10'b0000110100;
    parameter RCV_TERM_GND = "FALSE";
    parameter RCV_TERM_VTTRX = "TRUE";
    parameter RXGEARBOX_USE = "FALSE";
    parameter [23:0] RXPLL_COM_CFG = 24'h21680A;
    parameter [7:0] RXPLL_CP_CFG = 8'h00;
    parameter integer RXPLL_DIVSEL45_FB = 5;
    parameter integer RXPLL_DIVSEL_FB = 2;
    parameter integer RXPLL_DIVSEL_OUT = 1;
    parameter integer RXPLL_DIVSEL_REF = 1;
    parameter [2:0] RXPLL_LKDET_CFG = 3'b111;
    parameter [0:0] RXPRBSERR_LOOPBACK = 1'b0;
    parameter RXRECCLK_CTRL = "RXRECCLKPCS";
    parameter [9:0] RXRECCLK_DLY = 10'b0000000000;
    parameter [15:0] RXUSRCLK_DLY = 16'h0000;
    parameter RX_BUFFER_USE = "TRUE";
    parameter integer RX_CLK25_DIVIDER = 6;
    parameter integer RX_DATA_WIDTH = 20;
    parameter RX_DECODE_SEQ_MATCH = "TRUE";
    parameter [3:0] RX_DLYALIGN_CTRINC = 4'b0100;
    parameter [4:0] RX_DLYALIGN_EDGESET = 5'b00110;
    parameter [3:0] RX_DLYALIGN_LPFINC = 4'b0111;
    parameter [2:0] RX_DLYALIGN_MONSEL = 3'b000;
    parameter [7:0] RX_DLYALIGN_OVRDSETTING = 8'b00000000;
    parameter RX_EN_IDLE_HOLD_CDR = "FALSE";
    parameter RX_EN_IDLE_HOLD_DFE = "TRUE";
    parameter RX_EN_IDLE_RESET_BUF = "TRUE";
    parameter RX_EN_IDLE_RESET_FR = "TRUE";
    parameter RX_EN_IDLE_RESET_PH = "TRUE";
    parameter RX_EN_MODE_RESET_BUF = "TRUE";
    parameter RX_EN_RATE_RESET_BUF = "TRUE";
    parameter RX_EN_REALIGN_RESET_BUF = "FALSE";
    parameter RX_EN_REALIGN_RESET_BUF2 = "FALSE";
    parameter [7:0] RX_EYE_OFFSET = 8'h4C;
    parameter [1:0] RX_EYE_SCANMODE = 2'b00;
    parameter RX_FIFO_ADDR_MODE = "FULL";
    parameter [3:0] RX_IDLE_HI_CNT = 4'b1000;
    parameter [3:0] RX_IDLE_LO_CNT = 4'b0000;
    parameter RX_LOSS_OF_SYNC_FSM = "FALSE";
    parameter integer RX_LOS_INVALID_INCR = 1;
    parameter integer RX_LOS_THRESHOLD = 4;
    parameter RX_OVERSAMPLE_MODE = "FALSE";
    parameter integer RX_SLIDE_AUTO_WAIT = 5;
    parameter RX_SLIDE_MODE = "OFF";
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COMSAS = 52;
    parameter integer SAS_MIN_COMSAS = 40;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter [2:0] SATA_IDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 7;
    parameter integer SATA_MAX_INIT = 22;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter integer SIM_GTXRESET_SPEEDUP = 1;
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter [2:0] SIM_RXREFCLK_SOURCE = 3'b000;
    parameter [2:0] SIM_TXREFCLK_SOURCE = 3'b000;
    parameter SIM_TX_ELEC_IDLE_LEVEL = "X";
    parameter SIM_VERSION = "2.0";
    parameter [4:0] TERMINATION_CTRL = 5'b10100;
    parameter TERMINATION_OVRD = "FALSE";
    parameter [11:0] TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] TRANS_TIME_NON_P2 = 8'h19;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [9:0] TRANS_TIME_TO_P2 = 10'h064;
    parameter [31:0] TST_ATTR = 32'h00000000;
    parameter TXDRIVE_LOOPBACK_HIZ = "FALSE";
    parameter TXDRIVE_LOOPBACK_PD = "FALSE";
    parameter TXGEARBOX_USE = "FALSE";
    parameter TXOUTCLK_CTRL = "TXOUTCLKPCS";
    parameter [9:0] TXOUTCLK_DLY = 10'b0000000000;
    parameter [23:0] TXPLL_COM_CFG = 24'h21680A;
    parameter [7:0] TXPLL_CP_CFG = 8'h00;
    parameter integer TXPLL_DIVSEL45_FB = 5;
    parameter integer TXPLL_DIVSEL_FB = 2;
    parameter integer TXPLL_DIVSEL_OUT = 1;
    parameter integer TXPLL_DIVSEL_REF = 1;
    parameter [2:0] TXPLL_LKDET_CFG = 3'b111;
    parameter [1:0] TXPLL_SATA = 2'b00;
    parameter TX_BUFFER_USE = "TRUE";
    parameter [5:0] TX_BYTECLK_CFG = 6'h00;
    parameter integer TX_CLK25_DIVIDER = 6;
    parameter TX_CLK_SOURCE = "RXPLL";
    parameter integer TX_DATA_WIDTH = 20;
    parameter [4:0] TX_DEEMPH_0 = 5'b11010;
    parameter [4:0] TX_DEEMPH_1 = 5'b10000;
    parameter [13:0] TX_DETECT_RX_CFG = 14'h1832;
    parameter [3:0] TX_DLYALIGN_CTRINC = 4'b0100;
    parameter [3:0] TX_DLYALIGN_LPFINC = 4'b0110;
    parameter [2:0] TX_DLYALIGN_MONSEL = 3'b000;
    parameter [7:0] TX_DLYALIGN_OVRDSETTING = 8'b10000000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter TX_EN_RATE_RESET_BUF = "TRUE";
    parameter [2:0] TX_IDLE_ASSERT_DELAY = 3'b100;
    parameter [2:0] TX_IDLE_DEASSERT_DELAY = 3'b010;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter TX_OVERSAMPLE_MODE = "FALSE";
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [1:0] TX_TDCC_CFG = 2'b11;
    parameter [5:0] TX_USRCLK_CFG = 6'h00;
    parameter TX_XCLK_SEL = "TXUSR";
    output COMFINISH;
    output COMINITDET;
    output COMSASDET;
    output COMWAKEDET;
    output DRDY;
    output PHYSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMMADET;
    output RXDATAVALID;
    output RXELECIDLE;
    output RXHEADERVALID;
    output RXOVERSAMPLEERR;
    output RXPLLLKDET;
    output RXPRBSERR;
    output RXRATEDONE;
    output RXRECCLK;
    output RXRECCLKPCS;
    output RXRESETDONE;
    output RXSTARTOFSEQ;
    output RXVALID;
    output TXGEARBOXREADY;
    output TXN;
    output TXOUTCLK;
    output TXOUTCLKPCS;
    output TXP;
    output TXPLLLKDET;
    output TXRATEDONE;
    output TXRESETDONE;
    output [15:0] DRPDO;
    output [1:0] MGTREFCLKFAB;
    output [1:0] RXLOSSOFSYNC;
    output [1:0] TXBUFSTATUS;
    output [2:0] DFESENSCAL;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXCLKCORCNT;
    output [2:0] RXHEADER;
    output [2:0] RXSTATUS;
    output [31:0] RXDATA;
    output [3:0] DFETAP3MONITOR;
    output [3:0] DFETAP4MONITOR;
    output [3:0] RXCHARISCOMMA;
    output [3:0] RXCHARISK;
    output [3:0] RXCHBONDO;
    output [3:0] RXDISPERR;
    output [3:0] RXNOTINTABLE;
    output [3:0] RXRUNDISP;
    output [3:0] TXKERR;
    output [3:0] TXRUNDISP;
    output [4:0] DFEEYEDACMON;
    output [4:0] DFETAP1MONITOR;
    output [4:0] DFETAP2MONITOR;
    output [5:0] DFECLKDLYADJMON;
    output [7:0] RXDLYALIGNMONITOR;
    output [7:0] TXDLYALIGNMONITOR;
    output [9:0] TSTOUT;
    input DCLK;
    input DEN;
    input DFEDLYOVRD;
    input DFETAPOVRD;
    input DWE;
    input GATERXELECIDLE;
    input GREFCLKRX;
    input GREFCLKTX;
    input GTXRXRESET;
    input GTXTXRESET;
    input IGNORESIGDET;
    input PERFCLKRX;
    input PERFCLKTX;
    input PLLRXRESET;
    input PLLTXRESET;
    input PRBSCNTRESET;
    input RXBUFRESET;
    input RXCDRRESET;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETUSE;
    input RXDEC8B10BUSE;
    input RXDLYALIGNDISABLE;
    input RXDLYALIGNMONENB;
    input RXDLYALIGNOVERRIDE;
    input RXDLYALIGNRESET;
    input RXDLYALIGNSWPPRECURB;
    input RXDLYALIGNUPDSW;
    input RXENCHANSYNC;
    input RXENMCOMMAALIGN;
    input RXENPCOMMAALIGN;
    input RXENPMAPHASEALIGN;
    input RXENSAMPLEALIGN;
    input RXGEARBOXSLIP;
    input RXN;
    input RXP;
    input RXPLLLKDETEN;
    input RXPLLPOWERDOWN;
    input RXPMASETPHASE;
    input RXPOLARITY;
    input RXRESET;
    input RXSLIDE;
    input RXUSRCLK2;
    input RXUSRCLK;
    input TSTCLK0;
    input TSTCLK1;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDLYALIGNDISABLE;
    input TXDLYALIGNMONENB;
    input TXDLYALIGNOVERRIDE;
    input TXDLYALIGNRESET;
    input TXDLYALIGNUPDSW;
    input TXELECIDLE;
    input TXENC8B10BUSE;
    input TXENPMAPHASEALIGN;
    input TXINHIBIT;
    input TXPDOWNASYNCH;
    input TXPLLLKDETEN;
    input TXPLLPOWERDOWN;
    input TXPMASETPHASE;
    input TXPOLARITY;
    input TXPRBSFORCEERR;
    input TXRESET;
    input TXSTARTSEQ;
    input TXSWING;
    input TXUSRCLK2;
    input TXUSRCLK;
    input USRCODEERR;
    input [12:0] GTXTEST;
    input [15:0] DI;
    input [19:0] TSTIN;
    input [1:0] MGTREFCLKRX;
    input [1:0] MGTREFCLKTX;
    input [1:0] NORTHREFCLKRX;
    input [1:0] NORTHREFCLKTX;
    input [1:0] RXPOWERDOWN;
    input [1:0] RXRATE;
    input [1:0] SOUTHREFCLKRX;
    input [1:0] SOUTHREFCLKTX;
    input [1:0] TXPOWERDOWN;
    input [1:0] TXRATE;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXENPRBSTST;
    input [2:0] RXPLLREFSELDY;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXENPRBSTST;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXPLLREFSELDY;
    input [31:0] TXDATA;
    input [3:0] DFETAP3;
    input [3:0] DFETAP4;
    input [3:0] RXCHBONDI;
    input [3:0] TXBYPASS8B10B;
    input [3:0] TXCHARDISPMODE;
    input [3:0] TXCHARDISPVAL;
    input [3:0] TXCHARISK;
    input [3:0] TXDIFFCTRL;
    input [3:0] TXPREEMPHASIS;
    input [4:0] DFETAP1;
    input [4:0] DFETAP2;
    input [4:0] TXPOSTEMPHASIS;
    input [5:0] DFECLKDLYADJ;
    input [6:0] TXSEQUENCE;
    input [7:0] DADDR;
    input [9:0] RXEQMIX;
endmodule

module IBUFDS_GTXE1 (...);
    parameter CLKCM_CFG = "TRUE";
    parameter CLKRCV_TRST = "TRUE";
    parameter [9:0] REFCLKOUT_DLY = 10'b0000000000;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_GTHE1 (...);
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module GTHE2_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [19:0] ADAPT_CFG0 = 20'h00C10;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [41:0] CFOK_CFG = 42'h24800040E80;
    parameter [5:0] CFOK_CFG2 = 6'b100000;
    parameter [5:0] CFOK_CFG3 = 6'b100000;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 1;
    parameter [28:0] CPLL_CFG = 29'h00BC07DC;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 5;
    parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [23:0] DMONITOR_CFG = 24'h000A00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "TRUE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
    parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
    parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
    parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [2:0] GEARBOX_MODE = 3'b000;
    parameter [0:0] IS_CLKRSVD0_INVERTED = 1'b0;
    parameter [0:0] IS_CLKRSVD1_INVERTED = 1'b0;
    parameter [0:0] IS_CPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DMONITORCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_SIGVALIDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXPHDLYTSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] LOOPBACK_CFG = 1'b0;
    parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [31:0] PMA_RSV = 32'b00000000000000000000000010000000;
    parameter [31:0] PMA_RSV2 = 32'b00011100000000000000000000001010;
    parameter [1:0] PMA_RSV3 = 2'b00;
    parameter [14:0] PMA_RSV4 = 15'b000000000001000;
    parameter [3:0] PMA_RSV5 = 4'b0000;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 61;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [82:0] RXCDR_CFG = 83'h0002007FE2000C208001A;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [8:0] RXDLY_LCFG = 9'h030;
    parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [13:0] RXLPM_HF_CFG = 14'b00001000000000;
    parameter [17:0] RXLPM_LF_CFG = 18'b001001000000000000;
    parameter [6:0] RXOOB_CFG = 7'b0000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter [4:0] RXOSCALRESET_TIMEOUT = 5'b00000;
    parameter integer RXOUT_DIV = 2;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [23:0] RXPHDLY_CFG = 24'h084020;
    parameter [23:0] RXPH_CFG = 24'hC00002;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] RXPI_CFG0 = 2'b00;
    parameter [1:0] RXPI_CFG1 = 2'b00;
    parameter [1:0] RXPI_CFG2 = 2'b00;
    parameter [1:0] RXPI_CFG3 = 2'b00;
    parameter [0:0] RXPI_CFG4 = 1'b0;
    parameter [0:0] RXPI_CFG5 = 1'b0;
    parameter [2:0] RXPI_CFG6 = 3'b100;
    parameter [4:0] RXPMARESET_TIME = 5'b00011;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [23:0] RX_BIAS_CFG = 24'b000011000000000000010000;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter integer RX_CLK25_DIV = 7;
    parameter [0:0] RX_CLKMUX_PD = 1'b1;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter [13:0] RX_DEBUG_CFG = 14'b00000000000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [3:0] RX_DFELPM_CFG0 = 4'b0110;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter [2:0] RX_DFE_AGC_CFG1 = 3'b010;
    parameter [3:0] RX_DFE_AGC_CFG2 = 4'b0000;
    parameter [0:0] RX_DFE_AGC_OVRDEN = 1'b1;
    parameter [22:0] RX_DFE_GAIN_CFG = 23'h0020C0;
    parameter [11:0] RX_DFE_H2_CFG = 12'b000000000000;
    parameter [11:0] RX_DFE_H3_CFG = 12'b000001000000;
    parameter [10:0] RX_DFE_H4_CFG = 11'b00011100000;
    parameter [10:0] RX_DFE_H5_CFG = 11'b00011100000;
    parameter [10:0] RX_DFE_H6_CFG = 11'b00000100000;
    parameter [10:0] RX_DFE_H7_CFG = 11'b00000100000;
    parameter [32:0] RX_DFE_KL_CFG = 33'b000000000000000000000001100010000;
    parameter [1:0] RX_DFE_KL_LPM_KH_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KH_CFG1 = 3'b010;
    parameter [3:0] RX_DFE_KL_LPM_KH_CFG2 = 4'b0010;
    parameter [0:0] RX_DFE_KL_LPM_KH_OVRDEN = 1'b1;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b10;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [3:0] RX_DFE_KL_LPM_KL_CFG2 = 4'b0010;
    parameter [0:0] RX_DFE_KL_LPM_KL_OVRDEN = 1'b1;
    parameter [15:0] RX_DFE_LPM_CFG = 16'h0080;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter [53:0] RX_DFE_ST_CFG = 54'h00E100000C003F;
    parameter [16:0] RX_DFE_UT_CFG = 17'b00011100000000000;
    parameter [16:0] RX_DFE_VP_CFG = 17'b00011101010100011;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter integer RX_INT_DATAWIDTH = 0;
    parameter [12:0] RX_OS_CFG = 13'b0000010000000;
    parameter integer RX_SIG_VALID_DLY = 10;
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
    parameter SIM_VERSION = "1.1";
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [31:0] TST_RSV = 32'h00000000;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [8:0] TXDLY_LCFG = 9'h030;
    parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
    parameter TXGEARBOX_EN = "FALSE";
    parameter [0:0] TXOOB_CFG = 1'b0;
    parameter integer TXOUT_DIV = 2;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [23:0] TXPHDLY_CFG = 24'h084020;
    parameter [15:0] TXPH_CFG = 16'h0780;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b0;
    parameter [2:0] TXPI_CFG5 = 3'b100;
    parameter [0:0] TXPI_GREY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 7;
    parameter [0:0] TX_CLKMUX_PD = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter integer TX_INT_DATAWIDTH = 0;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
    parameter [16:0] TX_RXDETECT_PRECHARGE_TIME = 17'h00000;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter TX_XCLK_SEL = "TXUSR";
    parameter [0:0] UCODEER_CLR = 1'b0;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTREFCLKMONITOR;
    output PHYSTATUS;
    output RSOSINTDONE;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output RXDFESLIDETAPSTARTED;
    output RXDFESLIDETAPSTROBEDONE;
    output RXDFESLIDETAPSTROBESTARTED;
    output RXDFESTADAPTDONE;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRESETDONE;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXGEARBOXREADY;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    output [14:0] DMONITOROUT;
    output [15:0] DRPDO;
    output [15:0] PCSRSVDOUT;
    output [1:0] RXCLKCORCNT;
    output [1:0] RXDATAVALID;
    output [1:0] RXHEADERVALID;
    output [1:0] RXSTARTOFSEQ;
    output [1:0] TXBUFSTATUS;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXSTATUS;
    output [4:0] RXCHBONDO;
    output [4:0] RXPHMONITOR;
    output [4:0] RXPHSLIPMONITOR;
    output [5:0] RXHEADER;
    output [63:0] RXDATA;
    output [6:0] RXMONITOROUT;
    output [7:0] RXCHARISCOMMA;
    output [7:0] RXCHARISK;
    output [7:0] RXDISPERR;
    output [7:0] RXNOTINTABLE;
    input CFGRESET;
    (* invertible_pin = "IS_CLKRSVD0_INVERTED" *)
    input CLKRSVD0;
    (* invertible_pin = "IS_CLKRSVD1_INVERTED" *)
    input CLKRSVD1;
    (* invertible_pin = "IS_CPLLLOCKDETCLK_INVERTED" *)
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input CPLLRESET;
    input DMONFIFORESET;
    (* invertible_pin = "IS_DMONITORCLK_INVERTED" *)
    input DMONITORCLK;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input QPLLCLK;
    input QPLLREFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input RXDDIEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFECM1EN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFESLIDETAPADAPTEN;
    input RXDFESLIDETAPHOLD;
    input RXDFESLIDETAPINITOVRDEN;
    input RXDFESLIDETAPONLYADAPTEN;
    input RXDFESLIDETAPOVRDEN;
    input RXDFESLIDETAPSTROBE;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input RXGEARBOXSLIP;
    input RXLPMEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXMCOMMAALIGNEN;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTNTRLEN;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input RXQPIEN;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input RXUSERRDY;
    (* invertible_pin = "IS_RXUSRCLK2_INVERTED" *)
    input RXUSRCLK2;
    (* invertible_pin = "IS_RXUSRCLK_INVERTED" *)
    input RXUSRCLK;
    input SETERRSTATUS;
    (* invertible_pin = "IS_SIGVALIDCLK_INVERTED" *)
    input SIGVALIDCLK;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXINHIBIT;
    input TXPCSRESET;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    (* invertible_pin = "IS_TXPHDLYTSTCLK_INVERTED" *)
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input TXPISOPD;
    input TXPMARESET;
    input TXPOLARITY;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input TXPRECURSORINV;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input TXRATEMODE;
    input TXSTARTSEQ;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input TXUSERRDY;
    (* invertible_pin = "IS_TXUSRCLK2_INVERTED" *)
    input TXUSRCLK2;
    (* invertible_pin = "IS_TXUSRCLK_INVERTED" *)
    input TXUSRCLK;
    input [13:0] RXADAPTSELTEST;
    input [15:0] DRPDI;
    input [15:0] GTRSVD;
    input [15:0] PCSRSVDIN;
    input [19:0] TSTIN;
    input [1:0] RXELECIDLEMODE;
    input [1:0] RXMONITORSEL;
    input [1:0] RXPD;
    input [1:0] RXSYSCLKSEL;
    input [1:0] TXPD;
    input [1:0] TXSYSCLKSEL;
    input [2:0] CPLLREFCLKSEL;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXOUTCLKSEL;
    input [2:0] RXPRBSSEL;
    input [2:0] RXRATE;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input [2:0] TXPRBSSEL;
    input [2:0] TXRATE;
    input [3:0] RXOSINTCFG;
    input [3:0] RXOSINTID0;
    input [3:0] TXDIFFCTRL;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input [4:0] RXCHBONDI;
    input [4:0] RXDFEAGCTRL;
    input [4:0] RXDFESLIDETAP;
    input [4:0] TXPIPPMSTEPSIZE;
    input [4:0] TXPOSTCURSOR;
    input [4:0] TXPRECURSOR;
    input [5:0] RXDFESLIDETAPID;
    input [63:0] TXDATA;
    input [6:0] TXMAINCURSOR;
    input [6:0] TXSEQUENCE;
    input [7:0] TX8B10BBYPASS;
    input [7:0] TXCHARDISPMODE;
    input [7:0] TXCHARDISPVAL;
    input [7:0] TXCHARISK;
    input [8:0] DRPADDR;
endmodule

module GTHE2_COMMON (...);
    parameter [63:0] BIAS_CFG = 64'h0000040000001000;
    parameter [31:0] COMMON_CFG = 32'h0000001C;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_QPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [26:0] QPLL_CFG = 27'h0480181;
    parameter [3:0] QPLL_CLKOUT_CFG = 4'b0000;
    parameter [5:0] QPLL_COARSE_FREQ_OVRD = 6'b010000;
    parameter [0:0] QPLL_COARSE_FREQ_OVRD_EN = 1'b0;
    parameter [9:0] QPLL_CP = 10'b0000011111;
    parameter [0:0] QPLL_CP_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_DMONITOR_SEL = 1'b0;
    parameter [9:0] QPLL_FBDIV = 10'b0000000000;
    parameter [0:0] QPLL_FBDIV_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_FBDIV_RATIO = 1'b0;
    parameter [23:0] QPLL_INIT_CFG = 24'h000006;
    parameter [15:0] QPLL_LOCK_CFG = 16'h01E8;
    parameter [3:0] QPLL_LPF = 4'b1111;
    parameter integer QPLL_REFCLK_DIV = 2;
    parameter [0:0] QPLL_RP_COMP = 1'b0;
    parameter [1:0] QPLL_VTRL_RESET = 2'b00;
    parameter [1:0] RCAL_CFG = 2'b00;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [2:0] SIM_QPLLREFCLK_SEL = 3'b001;
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_VERSION = "1.1";
    output DRPRDY;
    output QPLLFBCLKLOST;
    output QPLLLOCK;
    output QPLLOUTCLK;
    output QPLLOUTREFCLK;
    output QPLLREFCLKLOST;
    output REFCLKOUTMONITOR;
    output [15:0] DRPDO;
    output [15:0] PMARSVDOUT;
    output [7:0] QPLLDMONITOR;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input BGRCALOVRDENB;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    (* invertible_pin = "IS_QPLLLOCKDETCLK_INVERTED" *)
    input QPLLLOCKDETCLK;
    input QPLLLOCKEN;
    input QPLLOUTRESET;
    input QPLLPD;
    input QPLLRESET;
    input RCALENB;
    input [15:0] DRPDI;
    input [15:0] QPLLRSVD1;
    input [2:0] QPLLREFCLKSEL;
    input [4:0] BGRCALOVRD;
    input [4:0] QPLLRSVD2;
    input [7:0] DRPADDR;
    input [7:0] PMARSVD;
endmodule

module GTPE2_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [19:0] ADAPT_CFG0 = 20'b00000000000000000000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [42:0] CFOK_CFG = 43'b1001001000000000000000001000000111010000000;
    parameter [6:0] CFOK_CFG2 = 7'b0100000;
    parameter [6:0] CFOK_CFG3 = 7'b0100000;
    parameter [0:0] CFOK_CFG4 = 1'b0;
    parameter [1:0] CFOK_CFG5 = 2'b00;
    parameter [3:0] CFOK_CFG6 = 4'b0000;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter [0:0] CLK_COMMON_SWING = 1'b0;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 1;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [23:0] DMONITOR_CFG = 24'h000A00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h010;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
    parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
    parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
    parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [2:0] GEARBOX_MODE = 3'b000;
    parameter [0:0] IS_CLKRSVD0_INVERTED = 1'b0;
    parameter [0:0] IS_CLKRSVD1_INVERTED = 1'b0;
    parameter [0:0] IS_DMONITORCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_SIGVALIDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXPHDLYTSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] LOOPBACK_CFG = 1'b0;
    parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [0:0] PMA_LOOPBACK_CFG = 1'b0;
    parameter [31:0] PMA_RSV = 32'h00000333;
    parameter [31:0] PMA_RSV2 = 32'h00002050;
    parameter [1:0] PMA_RSV3 = 2'b00;
    parameter [3:0] PMA_RSV4 = 4'b0000;
    parameter [0:0] PMA_RSV5 = 1'b0;
    parameter [0:0] PMA_RSV6 = 1'b0;
    parameter [0:0] PMA_RSV7 = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 61;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [82:0] RXCDR_CFG = 83'h0000107FE406001041010;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [8:0] RXDLY_LCFG = 9'h020;
    parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [6:0] RXLPMRESET_TIME = 7'b0001111;
    parameter [0:0] RXLPM_BIAS_STARTUP_DISABLE = 1'b0;
    parameter [3:0] RXLPM_CFG = 4'b0110;
    parameter [0:0] RXLPM_CFG1 = 1'b0;
    parameter [0:0] RXLPM_CM_CFG = 1'b0;
    parameter [8:0] RXLPM_GC_CFG = 9'b111100010;
    parameter [2:0] RXLPM_GC_CFG2 = 3'b001;
    parameter [13:0] RXLPM_HF_CFG = 14'b00001111110000;
    parameter [4:0] RXLPM_HF_CFG2 = 5'b01010;
    parameter [3:0] RXLPM_HF_CFG3 = 4'b0000;
    parameter [0:0] RXLPM_HOLD_DURING_EIDLE = 1'b0;
    parameter [0:0] RXLPM_INCM_CFG = 1'b0;
    parameter [0:0] RXLPM_IPCM_CFG = 1'b0;
    parameter [17:0] RXLPM_LF_CFG = 18'b000000001111110000;
    parameter [4:0] RXLPM_LF_CFG2 = 5'b01010;
    parameter [2:0] RXLPM_OSINT_CFG = 3'b100;
    parameter [6:0] RXOOB_CFG = 7'b0000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter [4:0] RXOSCALRESET_TIMEOUT = 5'b00000;
    parameter integer RXOUT_DIV = 2;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [23:0] RXPHDLY_CFG = 24'h084000;
    parameter [23:0] RXPH_CFG = 24'hC00002;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [2:0] RXPI_CFG0 = 3'b000;
    parameter [0:0] RXPI_CFG1 = 1'b0;
    parameter [0:0] RXPI_CFG2 = 1'b0;
    parameter [4:0] RXPMARESET_TIME = 5'b00011;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [15:0] RX_BIAS_CFG = 16'b0000111100110011;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter integer RX_CLK25_DIV = 7;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter [13:0] RX_DEBUG_CFG = 14'b00000000000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [12:0] RX_OS_CFG = 13'b0001111110000;
    parameter integer RX_SIG_VALID_DLY = 10;
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SATA_PLL_CFG = "VCO_3000MHZ";
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
    parameter SIM_VERSION = "1.0";
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [31:0] TST_RSV = 32'h00000000;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [8:0] TXDLY_LCFG = 9'h020;
    parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
    parameter TXGEARBOX_EN = "FALSE";
    parameter [0:0] TXOOB_CFG = 1'b0;
    parameter integer TXOUT_DIV = 2;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [23:0] TXPHDLY_CFG = 24'h084000;
    parameter [15:0] TXPH_CFG = 16'h0400;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b0;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GREY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 7;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter TX_XCLK_SEL = "TXUSR";
    parameter [0:0] UCODEER_CLR = 1'b0;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPTXN;
    output GTPTXP;
    output PHYSTATUS;
    output PMARSVDOUT0;
    output PMARSVDOUT1;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output RXHEADERVALID;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXRATEDONE;
    output RXRESETDONE;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXGEARBOXREADY;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    output [14:0] DMONITOROUT;
    output [15:0] DRPDO;
    output [15:0] PCSRSVDOUT;
    output [1:0] RXCLKCORCNT;
    output [1:0] RXDATAVALID;
    output [1:0] RXSTARTOFSEQ;
    output [1:0] TXBUFSTATUS;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXHEADER;
    output [2:0] RXSTATUS;
    output [31:0] RXDATA;
    output [3:0] RXCHARISCOMMA;
    output [3:0] RXCHARISK;
    output [3:0] RXCHBONDO;
    output [3:0] RXDISPERR;
    output [3:0] RXNOTINTABLE;
    output [4:0] RXPHMONITOR;
    output [4:0] RXPHSLIPMONITOR;
    input CFGRESET;
    (* invertible_pin = "IS_CLKRSVD0_INVERTED" *)
    input CLKRSVD0;
    (* invertible_pin = "IS_CLKRSVD1_INVERTED" *)
    input CLKRSVD1;
    input DMONFIFORESET;
    (* invertible_pin = "IS_DMONITORCLK_INVERTED" *)
    input DMONITORCLK;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTPRXN;
    input GTPRXP;
    input GTRESETSEL;
    input GTRXRESET;
    input GTTXRESET;
    input PLL0CLK;
    input PLL0REFCLK;
    input PLL1CLK;
    input PLL1REFCLK;
    input PMARSVDIN0;
    input PMARSVDIN1;
    input PMARSVDIN2;
    input PMARSVDIN3;
    input PMARSVDIN4;
    input RESETOVRD;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input RXDDIEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input RXGEARBOXSLIP;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFOVRDEN;
    input RXLPMOSINTNTRLEN;
    input RXLPMRESET;
    input RXMCOMMAALIGNEN;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTNTRLEN;
    input RXOSINTOVRDEN;
    input RXOSINTPD;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input RXUSERRDY;
    (* invertible_pin = "IS_RXUSRCLK2_INVERTED" *)
    input RXUSRCLK2;
    (* invertible_pin = "IS_RXUSRCLK_INVERTED" *)
    input RXUSRCLK;
    input SETERRSTATUS;
    (* invertible_pin = "IS_SIGVALIDCLK_INVERTED" *)
    input SIGVALIDCLK;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXINHIBIT;
    input TXPCSRESET;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    (* invertible_pin = "IS_TXPHDLYTSTCLK_INVERTED" *)
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input TXPISOPD;
    input TXPMARESET;
    input TXPOLARITY;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input TXPRECURSORINV;
    input TXRATEMODE;
    input TXSTARTSEQ;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input TXUSERRDY;
    (* invertible_pin = "IS_TXUSRCLK2_INVERTED" *)
    input TXUSRCLK2;
    (* invertible_pin = "IS_TXUSRCLK_INVERTED" *)
    input TXUSRCLK;
    input [13:0] RXADAPTSELTEST;
    input [15:0] DRPDI;
    input [15:0] GTRSVD;
    input [15:0] PCSRSVDIN;
    input [19:0] TSTIN;
    input [1:0] RXELECIDLEMODE;
    input [1:0] RXPD;
    input [1:0] RXSYSCLKSEL;
    input [1:0] TXPD;
    input [1:0] TXSYSCLKSEL;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXOUTCLKSEL;
    input [2:0] RXPRBSSEL;
    input [2:0] RXRATE;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input [2:0] TXPRBSSEL;
    input [2:0] TXRATE;
    input [31:0] TXDATA;
    input [3:0] RXCHBONDI;
    input [3:0] RXOSINTCFG;
    input [3:0] RXOSINTID0;
    input [3:0] TX8B10BBYPASS;
    input [3:0] TXCHARDISPMODE;
    input [3:0] TXCHARDISPVAL;
    input [3:0] TXCHARISK;
    input [3:0] TXDIFFCTRL;
    input [4:0] TXPIPPMSTEPSIZE;
    input [4:0] TXPOSTCURSOR;
    input [4:0] TXPRECURSOR;
    input [6:0] TXMAINCURSOR;
    input [6:0] TXSEQUENCE;
    input [8:0] DRPADDR;
endmodule

module GTPE2_COMMON (...);
    parameter [63:0] BIAS_CFG = 64'h0000000000000000;
    parameter [31:0] COMMON_CFG = 32'h00000000;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK0_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK1_INVERTED = 1'b0;
    parameter [0:0] IS_PLL0LOCKDETCLK_INVERTED = 1'b0;
    parameter [0:0] IS_PLL1LOCKDETCLK_INVERTED = 1'b0;
    parameter [26:0] PLL0_CFG = 27'h01F03DC;
    parameter [0:0] PLL0_DMON_CFG = 1'b0;
    parameter integer PLL0_FBDIV = 4;
    parameter integer PLL0_FBDIV_45 = 5;
    parameter [23:0] PLL0_INIT_CFG = 24'h00001E;
    parameter [8:0] PLL0_LOCK_CFG = 9'h1E8;
    parameter integer PLL0_REFCLK_DIV = 1;
    parameter [26:0] PLL1_CFG = 27'h01F03DC;
    parameter [0:0] PLL1_DMON_CFG = 1'b0;
    parameter integer PLL1_FBDIV = 4;
    parameter integer PLL1_FBDIV_45 = 5;
    parameter [23:0] PLL1_INIT_CFG = 24'h00001E;
    parameter [8:0] PLL1_LOCK_CFG = 9'h1E8;
    parameter integer PLL1_REFCLK_DIV = 1;
    parameter [7:0] PLL_CLKOUT_CFG = 8'b00000000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [2:0] SIM_PLL0REFCLK_SEL = 3'b001;
    parameter [2:0] SIM_PLL1REFCLK_SEL = 3'b001;
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_VERSION = "1.0";
    output DRPRDY;
    output PLL0FBCLKLOST;
    output PLL0LOCK;
    output PLL0OUTCLK;
    output PLL0OUTREFCLK;
    output PLL0REFCLKLOST;
    output PLL1FBCLKLOST;
    output PLL1LOCK;
    output PLL1OUTCLK;
    output PLL1OUTREFCLK;
    output PLL1REFCLKLOST;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [15:0] DRPDO;
    output [15:0] PMARSVDOUT;
    output [7:0] DMONITOROUT;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input BGRCALOVRDENB;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input GTEASTREFCLK0;
    input GTEASTREFCLK1;
    (* invertible_pin = "IS_GTGREFCLK0_INVERTED" *)
    input GTGREFCLK0;
    (* invertible_pin = "IS_GTGREFCLK1_INVERTED" *)
    input GTGREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTWESTREFCLK0;
    input GTWESTREFCLK1;
    (* invertible_pin = "IS_PLL0LOCKDETCLK_INVERTED" *)
    input PLL0LOCKDETCLK;
    input PLL0LOCKEN;
    input PLL0PD;
    input PLL0RESET;
    (* invertible_pin = "IS_PLL1LOCKDETCLK_INVERTED" *)
    input PLL1LOCKDETCLK;
    input PLL1LOCKEN;
    input PLL1PD;
    input PLL1RESET;
    input RCALENB;
    input [15:0] DRPDI;
    input [15:0] PLLRSVD1;
    input [2:0] PLL0REFCLKSEL;
    input [2:0] PLL1REFCLKSEL;
    input [4:0] BGRCALOVRD;
    input [4:0] PLLRSVD2;
    input [7:0] DRPADDR;
    input [7:0] PMARSVD;
endmodule

module GTXE2_CHANNEL (...);
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 1;
    parameter [23:0] CPLL_CFG = 24'hB007D8;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 5;
    parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [23:0] DMONITOR_CFG = 24'h000A00;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
    parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
    parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
    parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [2:0] GEARBOX_MODE = 3'b000;
    parameter [0:0] IS_CPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXPHDLYTSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK_INVERTED = 1'b0;
    parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [31:0] PMA_RSV = 32'h00000000;
    parameter [15:0] PMA_RSV2 = 16'h2050;
    parameter [1:0] PMA_RSV3 = 2'b00;
    parameter [31:0] PMA_RSV4 = 32'h00000000;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 61;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [71:0] RXCDR_CFG = 72'h0B000023FF20400020;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [5:0] RXCDR_LOCK_CFG = 6'b010101;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [8:0] RXDLY_LCFG = 9'h030;
    parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [13:0] RXLPM_HF_CFG = 14'b00000011110000;
    parameter [13:0] RXLPM_LF_CFG = 14'b00000011110000;
    parameter [6:0] RXOOB_CFG = 7'b0000110;
    parameter integer RXOUT_DIV = 2;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [23:0] RXPHDLY_CFG = 24'h084020;
    parameter [23:0] RXPH_CFG = 24'h000000;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [4:0] RXPMARESET_TIME = 5'b00011;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [11:0] RX_BIAS_CFG = 12'b000000000000;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter integer RX_CLK25_DIV = 7;
    parameter [0:0] RX_CLKMUX_PD = 1'b1;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [2:0] RX_CM_TRIM = 3'b100;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter [11:0] RX_DEBUG_CFG = 12'b000000000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [22:0] RX_DFE_GAIN_CFG = 23'h180E0F;
    parameter [11:0] RX_DFE_H2_CFG = 12'b000111100000;
    parameter [11:0] RX_DFE_H3_CFG = 12'b000111100000;
    parameter [10:0] RX_DFE_H4_CFG = 11'b00011110000;
    parameter [10:0] RX_DFE_H5_CFG = 11'b00011110000;
    parameter [12:0] RX_DFE_KL_CFG = 13'b0001111110000;
    parameter [31:0] RX_DFE_KL_CFG2 = 32'h3008E56A;
    parameter [15:0] RX_DFE_LPM_CFG = 16'h0904;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter [16:0] RX_DFE_UT_CFG = 17'b00111111000000000;
    parameter [16:0] RX_DFE_VP_CFG = 17'b00011111100000000;
    parameter [12:0] RX_DFE_XYD_CFG = 13'b0000000010000;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter integer RX_INT_DATAWIDTH = 0;
    parameter [12:0] RX_OS_CFG = 13'b0001111110000;
    parameter integer RX_SIG_VALID_DLY = 10;
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
    parameter SIM_VERSION = "4.0";
    parameter [4:0] TERM_RCAL_CFG = 5'b10000;
    parameter [0:0] TERM_RCAL_OVRD = 1'b0;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [31:0] TST_RSV = 32'h00000000;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [8:0] TXDLY_LCFG = 9'h030;
    parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 2;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [23:0] TXPHDLY_CFG = 24'h084020;
    parameter [15:0] TXPH_CFG = 16'h0780;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter integer TX_CLK25_DIV = 7;
    parameter [0:0] TX_CLKMUX_PD = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [4:0] TX_DEEMPH0 = 5'b00000;
    parameter [4:0] TX_DEEMPH1 = 5'b00000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter integer TX_INT_DATAWIDTH = 0;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter TX_XCLK_SEL = "TXUSR";
    parameter [0:0] UCODEER_CLR = 1'b0;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTREFCLKMONITOR;
    output GTXTXN;
    output GTXTXP;
    output PHYSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output RXHEADERVALID;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPRBSERR;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRESETDONE;
    output RXSTARTOFSEQ;
    output RXVALID;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXGEARBOXREADY;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output [15:0] DRPDO;
    output [15:0] PCSRSVDOUT;
    output [1:0] RXCLKCORCNT;
    output [1:0] TXBUFSTATUS;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXHEADER;
    output [2:0] RXSTATUS;
    output [4:0] RXCHBONDO;
    output [4:0] RXPHMONITOR;
    output [4:0] RXPHSLIPMONITOR;
    output [63:0] RXDATA;
    output [6:0] RXMONITOROUT;
    output [7:0] DMONITOROUT;
    output [7:0] RXCHARISCOMMA;
    output [7:0] RXCHARISK;
    output [7:0] RXDISPERR;
    output [7:0] RXNOTINTABLE;
    output [9:0] TSTOUT;
    input CFGRESET;
    (* invertible_pin = "IS_CPLLLOCKDETCLK_INVERTED" *)
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input CPLLRESET;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTXRXN;
    input GTXRXP;
    input QPLLCLK;
    input QPLLREFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input RXDDIEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFECM1EN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDFEXYDHOLD;
    input RXDFEXYDOVRDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input RXGEARBOXSLIP;
    input RXLPMEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXMCOMMAALIGNEN;
    input RXOOBRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input RXQPIEN;
    input RXSLIDE;
    input RXUSERRDY;
    (* invertible_pin = "IS_RXUSRCLK2_INVERTED" *)
    input RXUSRCLK2;
    (* invertible_pin = "IS_RXUSRCLK_INVERTED" *)
    input RXUSRCLK;
    input SETERRSTATUS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXINHIBIT;
    input TXPCSRESET;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    (* invertible_pin = "IS_TXPHDLYTSTCLK_INVERTED" *)
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPISOPD;
    input TXPMARESET;
    input TXPOLARITY;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input TXPRECURSORINV;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input TXSTARTSEQ;
    input TXSWING;
    input TXUSERRDY;
    (* invertible_pin = "IS_TXUSRCLK2_INVERTED" *)
    input TXUSRCLK2;
    (* invertible_pin = "IS_TXUSRCLK_INVERTED" *)
    input TXUSRCLK;
    input [15:0] DRPDI;
    input [15:0] GTRSVD;
    input [15:0] PCSRSVDIN;
    input [19:0] TSTIN;
    input [1:0] RXELECIDLEMODE;
    input [1:0] RXMONITORSEL;
    input [1:0] RXPD;
    input [1:0] RXSYSCLKSEL;
    input [1:0] TXPD;
    input [1:0] TXSYSCLKSEL;
    input [2:0] CPLLREFCLKSEL;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXOUTCLKSEL;
    input [2:0] RXPRBSSEL;
    input [2:0] RXRATE;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input [2:0] TXPRBSSEL;
    input [2:0] TXRATE;
    input [3:0] CLKRSVD;
    input [3:0] TXDIFFCTRL;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN2;
    input [4:0] PMARSVDIN;
    input [4:0] RXCHBONDI;
    input [4:0] TXPOSTCURSOR;
    input [4:0] TXPRECURSOR;
    input [63:0] TXDATA;
    input [6:0] TXMAINCURSOR;
    input [6:0] TXSEQUENCE;
    input [7:0] TX8B10BBYPASS;
    input [7:0] TXCHARDISPMODE;
    input [7:0] TXCHARDISPVAL;
    input [7:0] TXCHARISK;
    input [8:0] DRPADDR;
endmodule

module GTXE2_COMMON (...);
    parameter [63:0] BIAS_CFG = 64'h0000040000001000;
    parameter [31:0] COMMON_CFG = 32'h00000000;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_QPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [26:0] QPLL_CFG = 27'h0680181;
    parameter [3:0] QPLL_CLKOUT_CFG = 4'b0000;
    parameter [5:0] QPLL_COARSE_FREQ_OVRD = 6'b010000;
    parameter [0:0] QPLL_COARSE_FREQ_OVRD_EN = 1'b0;
    parameter [9:0] QPLL_CP = 10'b0000011111;
    parameter [0:0] QPLL_CP_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_DMONITOR_SEL = 1'b0;
    parameter [9:0] QPLL_FBDIV = 10'b0000000000;
    parameter [0:0] QPLL_FBDIV_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_FBDIV_RATIO = 1'b0;
    parameter [23:0] QPLL_INIT_CFG = 24'h000006;
    parameter [15:0] QPLL_LOCK_CFG = 16'h21E8;
    parameter [3:0] QPLL_LPF = 4'b1111;
    parameter integer QPLL_REFCLK_DIV = 2;
    parameter [2:0] SIM_QPLLREFCLK_SEL = 3'b001;
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_VERSION = "4.0";
    output DRPRDY;
    output QPLLFBCLKLOST;
    output QPLLLOCK;
    output QPLLOUTCLK;
    output QPLLOUTREFCLK;
    output QPLLREFCLKLOST;
    output REFCLKOUTMONITOR;
    output [15:0] DRPDO;
    output [7:0] QPLLDMONITOR;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    (* invertible_pin = "IS_QPLLLOCKDETCLK_INVERTED" *)
    input QPLLLOCKDETCLK;
    input QPLLLOCKEN;
    input QPLLOUTRESET;
    input QPLLPD;
    input QPLLRESET;
    input RCALENB;
    input [15:0] DRPDI;
    input [15:0] QPLLRSVD1;
    input [2:0] QPLLREFCLKSEL;
    input [4:0] BGRCALOVRD;
    input [4:0] QPLLRSVD2;
    input [7:0] DRPADDR;
    input [7:0] PMARSVD;
endmodule

module IBUFDS_GTE2 (...);
    parameter CLKCM_CFG = "TRUE";
    parameter CLKRCV_TRST = "TRUE";
    parameter CLKSWING_CFG = "TRUE";
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module GTHE3_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'hF800;
    parameter [15:0] ADAPT_CFG1 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h20F8;
    parameter [15:0] CPLL_CFG1 = 16'hA494;
    parameter [15:0] CPLL_CFG2 = 16'hF001;
    parameter [5:0] CPLL_CFG3 = 6'h00;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [7:0] CPLL_INIT_CFG1 = 8'h00;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DFE_D_X_REL_POS = 1'b0;
    parameter [0:0] DFE_VCM_COMP_EN = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [10:0] EVODD_PHI_CFG = 11'b00000000000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] GM_BIAS_SELECT = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [2:0] PCS_RSVD1 = 3'b000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [1:0] PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [15:0] PMA_RSV1 = 16'h0000;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0000;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG1 = 16'h0080;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h07E6;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG4 = 16'h0000;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG5 = 16'h0000;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h0000;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h5080;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h07E0;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h7C42;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h4000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0060;
    parameter [15:0] RXCFOK_CFG2 = 16'h000E;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0032;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_CFG0 = 16'h0A00;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h7840;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h8000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h8000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_VP_CFG0 = 16'hAA00;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0033;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "Sigcfg_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h8000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0002;
    parameter [8:0] RXOOB_CFG = 9'b000000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h6622;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] RXPI_CFG0 = 2'b00;
    parameter [1:0] RXPI_CFG1 = 2'b00;
    parameter [1:0] RXPI_CFG2 = 2'b00;
    parameter [1:0] RXPI_CFG3 = 2'b00;
    parameter [0:0] RXPI_CFG4 = 1'b0;
    parameter [0:0] RXPI_CFG5 = 1'b1;
    parameter [2:0] RXPI_CFG6 = 3'b000;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h0AD4;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter [7:0] RX_CTLE3_LPF = 8'b00000000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [3:0] RX_DFELPM_CFG0 = 4'b0110;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter [2:0] RX_DFE_AGC_CFG1 = 3'b100;
    parameter [1:0] RX_DFE_KL_LPM_KH_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KH_CFG1 = 3'b010;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_HI_LR = 1'b0;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter real RX_PROGDIV_CFG = 4.0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter [1:0] RX_SUM_RES_CTRL = 2'b00;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b0000;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b000;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [0:0] RX_WIDEMODE_CDR = 1'b0;
    parameter RX_XCLK_SEL = "RXDES";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [0:0] SIM_TX_EIDLE_DRIVE_LEVEL = 1'b0;
    parameter integer SIM_VERSION = 2;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATUR_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter [3:0] TXDRVBIAS_N = 4'b1010;
    parameter [3:0] TXDRVBIAS_P = 4'b1100;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h2020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0001;
    parameter [15:0] TXPH_CFG = 16'h0980;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DCD_CFG = 6'b000010;
    parameter [0:0] TX_DCD_EN = 1'b0;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_EML_PHI_TUNE = 1'b0;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [2:0] TX_MODE_SEL = 3'b000;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 4.0;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [1:0] WB_MODE = 2'b00;
    output [2:0] BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output [2:0] BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [16:0] DMONITOROUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [11:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [7:0] PINRSRVDAS;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output [6:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [8:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input EVODDPHICALDONE;
    input EVODDPHICALSTART;
    input EVODDPHIDRDEN;
    input EVODDPHIDWREN;
    input EVODDPHIXRDEN;
    input EVODDPHIXWREN;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input [2:0] LOOPBACK;
    input LPBKRXTXSEREN;
    input LPBKTXRXSEREN;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input QPLL0CLK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RSTCLKENTX;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input [1:0] RXDFEAGCCTRL;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input [3:0] RXOSINTCFG;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input RXQPIEN;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input [2:0] TXBUFDIFFCTRL;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDEEMPH;
    input TXDETECTRX;
    input [3:0] TXDIFFCTRL;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPRECURSORINV;
    input TXPROGDIVRESET;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTHE3_COMMON (...);
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [9:0] BIAS_CFG_RSVD = 10'b0000000000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0004;
    parameter [15:0] QPLL0_CFG0 = 16'h3018;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0000;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0000;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0009;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h01E8;
    parameter [9:0] QPLL0_LPF = 10'b1111111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter integer QPLL0_REFCLK_DIV = 2;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'b0000000000000000;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] QPLL1_CFG0 = 16'h3018;
    parameter [15:0] QPLL1_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0000;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0000;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0009;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1111111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter integer QPLL1_REFCLK_DIV = 2;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'b0000000000000000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_EN = 1'b1;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0DATA1_0 = 16'b0000000000000000;
    parameter [8:0] SDM0DATA1_1 = 9'b000000000;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [0:0] SDM0_DATA_PIN_SEL = 1'b0;
    parameter [0:0] SDM0_WIDTH_PIN_SEL = 1'b0;
    parameter [15:0] SDM1DATA1_0 = 16'b0000000000000000;
    parameter [8:0] SDM1DATA1_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter [0:0] SDM1_DATA_PIN_SEL = 1'b0;
    parameter [0:0] SDM1_WIDTH_PIN_SEL = 1'b0;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer SIM_VERSION = 2;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0_SEL;
    output [1:0] RXRECCLK1_SEL;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [8:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
endmodule

module GTHE4_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_RXTERMINATION = 1'b1;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter [0:0] CAPBYPASS_FORCE = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter [0:0] CFOK_PWRSVE_EN = 1'b1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h2424;
    parameter [15:0] CKCAL1_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter [15:0] CKCAL_RSVD0 = 16'h4000;
    parameter [15:0] CKCAL_RSVD1 = 16'h0000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h01FA;
    parameter [15:0] CPLL_CFG1 = 16'h24A9;
    parameter [15:0] CPLL_CFG2 = 16'h6807;
    parameter [15:0] CPLL_CFG3 = 16'h0000;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DELAY_ELEC = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h800;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [2:0] LPBK_BIAS_CTRL = 3'b000;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter [2:0] LPBK_IND_CTRL0 = 3'b000;
    parameter [2:0] LPBK_IND_CTRL1 = 3'b000;
    parameter [2:0] LPBK_IND_CTRL2 = 3'b000;
    parameter [3:0] LPBK_RG_CTRL = 4'b0000;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'b00000;
    parameter [5:0] PCIE3_CLK_COR_FULL_THRSH = 6'b010000;
    parameter [4:0] PCIE3_CLK_COR_MAX_LAT = 5'b01000;
    parameter [4:0] PCIE3_CLK_COR_MIN_LAT = 5'b00100;
    parameter [5:0] PCIE3_CLK_COR_THRSH_TIMER = 6'b001000;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN4 = 2'h0;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0;
    parameter [0:0] RCLK_SIPO_INV_EN = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [2:0] RTX_BUF_CML_CTRL = 3'b010;
    parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0003;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0003;
    parameter [15:0] RXCDR_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h0164;
    parameter [9:0] RXCDR_CFG2_GEN2 = 10'h164;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0034;
    parameter [15:0] RXCDR_CFG2_GEN4 = 16'h0034;
    parameter [15:0] RXCDR_CFG3 = 16'h0024;
    parameter [5:0] RXCDR_CFG3_GEN2 = 6'h24;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0024;
    parameter [15:0] RXCDR_CFG3_GEN4 = 16'h0024;
    parameter [15:0] RXCDR_CFG4 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG5 = 16'hB46B;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h146B;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h0000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0002;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_KH_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG3 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0002;
    parameter [0:0] RXDFE_PWR_SAVING = 1'b0;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_UT_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h1000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000110000;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [0:0] RXPI_AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [15:0] RXPI_CFG0 = 16'h0002;
    parameter [15:0] RXPI_CFG1 = 16'b0000000000000000;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [1:0] RXPI_SEL_LC = 2'b00;
    parameter [1:0] RXPI_STARTCODE = 2'b00;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter [0:0] RXREFCLKDIV2_SEL = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h12B0;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 12;
    parameter [7:0] RX_CTLE3_LPF = 8'b00000000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b011;
    parameter integer RX_DFELPM_CFG0 = 0;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b1;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 4;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [0:0] RX_DIV2_MODE_B = 1'b0;
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter [0:0] RX_EN_HI_LR = 1'b1;
    parameter [8:0] RX_EXT_RL_CTRL = 9'b000000000;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] RX_PMA_RSV0 = 16'h0000;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b1001;
    parameter [3:0] RX_SUM_RESLOAD_CTRL = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b1010;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b101;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter [0:0] SAMPLE_CLK_PHASE = 1'b0;
    parameter [0:0] SAS_12G_MODE = 1'b0;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
    parameter [0:0] SRSTMODE = 1'b0;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATURE_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter [3:0] TXDRVBIAS_N = 4'b1010;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h6020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0002;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] TXPI_CFG = 16'h0000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter [0:0] TXPI_PPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXREFCLKDIV2_SEL = 1'b0;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [5:0] TX_DEEMPH2 = 6'b000000;
    parameter [5:0] TX_DEEMPH3 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter integer TX_DRVMUX_CTRL = 2;
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h003F;
    parameter [15:0] TX_PHICAL_CFG2 = 16'h0000;
    parameter integer TX_PI_BIASSET = 0;
    parameter [1:0] TX_PI_IBIAS_MID = 2'b00;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] TX_PMA_RSV0 = 16'h0008;
    parameter integer TX_PREDRV_CTRL = 2;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 3;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter [1:0] TX_SW_MEAS = 2'b00;
    parameter [2:0] TX_VREG_CTRL = 3'b000;
    parameter [0:0] TX_VREG_PDB = 1'b0;
    parameter [1:0] TX_VREG_VREFSEL = 2'b00;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USB_BOTH_BURST_IDLE = 1'b0;
    parameter [6:0] USB_BURSTMAX_U3WAKE = 7'b1111111;
    parameter [6:0] USB_BURSTMIN_U3WAKE = 7'b1100011;
    parameter [0:0] USB_CLK_COR_EQ_EN = 1'b0;
    parameter [0:0] USB_EXT_CNTL = 1'b1;
    parameter [9:0] USB_IDLEMAX_POLLING = 10'b1010111011;
    parameter [9:0] USB_IDLEMIN_POLLING = 10'b0100101011;
    parameter [8:0] USB_LFPSPING_BURST = 9'b000000101;
    parameter [8:0] USB_LFPSPOLLING_BURST = 9'b000110001;
    parameter [8:0] USB_LFPSPOLLING_IDLE_MS = 9'b000000100;
    parameter [8:0] USB_LFPSU1EXIT_BURST = 9'b000011101;
    parameter [8:0] USB_LFPSU2LPEXIT_BURST_MS = 9'b001100011;
    parameter [8:0] USB_LFPSU3WAKE_BURST_MS = 9'b111110011;
    parameter [3:0] USB_LFPS_TPERIOD = 4'b0011;
    parameter [0:0] USB_LFPS_TPERIOD_ACCURATE = 1'b1;
    parameter [0:0] USB_MODE = 1'b0;
    parameter [0:0] USB_PCIE_ERR_REP_DIS = 1'b0;
    parameter integer USB_PING_SATA_MAX_INIT = 21;
    parameter integer USB_PING_SATA_MIN_INIT = 12;
    parameter integer USB_POLL_SATA_MAX_BURST = 8;
    parameter integer USB_POLL_SATA_MIN_BURST = 4;
    parameter [0:0] USB_RAW_ELEC = 1'b0;
    parameter [0:0] USB_RXIDLE_P0_CTRL = 1'b1;
    parameter [0:0] USB_TXIDLE_TUNE_ENABLE = 1'b1;
    parameter integer USB_U1_SATA_MAX_WAKE = 7;
    parameter integer USB_U1_SATA_MIN_WAKE = 4;
    parameter integer USB_U2_SAS_MAX_COM = 64;
    parameter integer USB_U2_SAS_MIN_COM = 36;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [0:0] Y_ALL_MODE = 1'b0;
    output BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [15:0] DMONITOROUT;
    output DMONITOROUTCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [15:0] PINRSRVDAS;
    output POWERPRESENT;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output RXLFPSTRESETDET;
    output RXLFPSU2LPEXITDET;
    output RXLFPSU3WAKEDET;
    output [7:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLFREQLOCK;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input FREQOS;
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTRXRESETSEL;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTTXRESETSEL;
    input INCPCTRL;
    input [2:0] LOOPBACK;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input QPLL0CLK;
    input QPLL0FREQLOCK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1FREQLOCK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXAFECFOKEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input [6:0] RXCKCALSTART;
    input RXCOMMADETEN;
    input [1:0] RXDFEAGCCTRL;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input [3:0] RXDFECFOKFCNUM;
    input RXDFECFOKFEN;
    input RXDFECFOKFPULSE;
    input RXDFECFOKHOLD;
    input RXDFECFOKOVREN;
    input RXDFEKHHOLD;
    input RXDFEKHOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXEQTRAINING;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input RXQPIEN;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXTERMINATION;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input [1:0] TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input TXLFPSTRESET;
    input TXLFPSU2LPEXIT;
    input TXLFPSU3WAKE;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input TXMUXDCDEXHOLD;
    input TXMUXDCDORWREN;
    input TXONESZEROS;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input TXQPIBIASEN;
    input TXQPIWEAKPUP;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTHE4_COMMON (...);
    parameter [0:0] AEN_QPLL0_FBDIV = 1'b1;
    parameter [0:0] AEN_QPLL1_FBDIV = 1'b1;
    parameter [0:0] AEN_SDM0TOGGLE = 1'b0;
    parameter [0:0] AEN_SDM1TOGGLE = 1'b0;
    parameter [0:0] A_SDM0TOGGLE = 1'b0;
    parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000;
    parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000;
    parameter [0:0] A_SDM1TOGGLE = 1'b0;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [15:0] BIAS_CFG_RSVD = 16'h0000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0000;
    parameter [15:0] PPF0_CFG = 16'h0F00;
    parameter [15:0] PPF1_CFG = 16'h0F00;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h391C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0F80;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0002;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1011111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL0_PCI_EN = 1'b0;
    parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL0_REFCLK_DIV = 1;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h691C;
    parameter [15:0] QPLL1_CFG1 = 16'h0020;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0F80;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0002;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1011111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL1_PCI_EN = 1'b0;
    parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL1_REFCLK_DIV = 1;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_ENB = 1'b0;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0SEL;
    output [1:0] RXRECCLK1SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    output [9:0] TCONGPO;
    output TCONRSVDOUT0;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [15:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [2:0] PCIERATEQPLL0;
    input [2:0] PCIERATEQPLL1;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input [7:0] QPLL0FBDIV;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input [7:0] QPLL1FBDIV;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input SDM0TOGGLE;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input SDM1TOGGLE;
    input [1:0] SDM1WIDTH;
    input [9:0] TCONGPI;
    input TCONPOWERUP;
    input [1:0] TCONRESET;
    input [1:0] TCONRSVDIN1;
endmodule

module GTYE3_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'b0000000000000000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter [0:0] CAPBYPASS_FORCE = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h0000;
    parameter [15:0] CKCAL1_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter [15:0] CKCAL_RSVD0 = 16'h0000;
    parameter [15:0] CKCAL_RSVD1 = 16'h0000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h20F8;
    parameter [15:0] CPLL_CFG1 = 16'hA494;
    parameter [15:0] CPLL_CFG2 = 16'hF001;
    parameter [5:0] CPLL_CFG3 = 6'h00;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [7:0] CPLL_INIT_CFG1 = 8'h00;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DFE_D_X_REL_POS = 1'b0;
    parameter [0:0] DFE_VCM_COMP_EN = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter [10:0] EVODD_PHI_CFG = 11'b00000000000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] GM_BIAS_SELECT = 1'b0;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [15:0] LOOP0_CFG = 16'h0000;
    parameter [15:0] LOOP10_CFG = 16'h0000;
    parameter [15:0] LOOP11_CFG = 16'h0000;
    parameter [15:0] LOOP12_CFG = 16'h0000;
    parameter [15:0] LOOP13_CFG = 16'h0000;
    parameter [15:0] LOOP1_CFG = 16'h0000;
    parameter [15:0] LOOP2_CFG = 16'h0000;
    parameter [15:0] LOOP3_CFG = 16'h0000;
    parameter [15:0] LOOP4_CFG = 16'h0000;
    parameter [15:0] LOOP5_CFG = 16'h0000;
    parameter [15:0] LOOP6_CFG = 16'h0000;
    parameter [15:0] LOOP7_CFG = 16'h0000;
    parameter [15:0] LOOP8_CFG = 16'h0000;
    parameter [15:0] LOOP9_CFG = 16'h0000;
    parameter [2:0] LPBK_BIAS_CTRL = 3'b000;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter [3:0] LPBK_RG_CTRL = 4'b0000;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [2:0] PCS_RSVD1 = 3'b000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [1:0] PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [15:0] PMA_RSV0 = 16'h0000;
    parameter [15:0] PMA_RSV1 = 16'h0000;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0000;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG1 = 16'h0300;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0300;
    parameter [15:0] RXCDR_CFG2 = 16'h0060;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0060;
    parameter [15:0] RXCDR_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG4 = 16'h0002;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h0002;
    parameter [15:0] RXCDR_CFG5 = 16'h0000;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h0000;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0001;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [1:0] RXCFOKDONE_SRC = 2'b00;
    parameter [15:0] RXCFOK_CFG0 = 16'h3E00;
    parameter [15:0] RXCFOK_CFG1 = 16'h0042;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4C00;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h1E00;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h1900;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0200;
    parameter [0:0] RXDFE_PWR_SAVING = 1'b0;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h0200;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0400;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [0:0] RXPI_AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [15:0] RXPI_CFG = 16'h0100;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [15:0] RXPI_RSV0 = 16'h0000;
    parameter [1:0] RXPI_SEL_LC = 2'b00;
    parameter [1:0] RXPI_STARTCODE = 2'b00;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h1534;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 10;
    parameter [0:0] RX_CTLE1_KHKL = 1'b0;
    parameter [0:0] RX_CTLE2_KHKL = 1'b0;
    parameter [0:0] RX_CTLE3_AGC = 1'b0;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b010;
    parameter integer RX_DFELPM_CFG0 = 6;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 2;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [0:0] RX_DIV2_MODE_B = 1'b0;
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter [0:0] RX_EN_HI_LR = 1'b0;
    parameter [8:0] RX_EXT_RL_CTRL = 9'b000000000;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b1000;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b101;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [0:0] SIM_TX_EIDLE_DRIVE_LEVEL = 1'b0;
    parameter integer SIM_VERSION = 2;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATURE_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h2020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0001;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [15:0] TXPI_RSV0 = 16'h0000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter [0:0] TX_CLKREG_PDB = 1'b0;
    parameter [2:0] TX_CLKREG_SET = 3'b000;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DCD_CFG = 6'b000010;
    parameter [0:0] TX_DCD_EN = 1'b0;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter integer TX_DRVMUX_CTRL = 2;
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_EML_PHI_TUNE = 1'b0;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [2:0] TX_MODE_SEL = 3'b000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h7E00;
    parameter [15:0] TX_PHICAL_CFG2 = 16'h0000;
    parameter integer TX_PI_BIASSET = 0;
    parameter [15:0] TX_PI_CFG0 = 16'h0000;
    parameter [15:0] TX_PI_CFG1 = 16'h0000;
    parameter [0:0] TX_PI_DIV2_MODE_B = 1'b0;
    parameter [0:0] TX_PI_SEL_QPLL0 = 1'b0;
    parameter [0:0] TX_PI_SEL_QPLL1 = 1'b0;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter integer TX_PREDRV_CTRL = 2;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 4;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output [2:0] BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output [2:0] BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [16:0] DMONITOROUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output GTYTXN;
    output GTYTXP;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [7:0] PINRSRVDAS;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output [6:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input ELPCALDVORWREN;
    input ELPCALPAORWREN;
    input EVODDPHICALDONE;
    input EVODDPHICALSTART;
    input EVODDPHIDRDEN;
    input EVODDPHIDWREN;
    input EVODDPHIXRDEN;
    input EVODDPHIXWREN;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTYRXN;
    input GTYRXP;
    input [2:0] LOOPBACK;
    input [15:0] LOOPRSVD;
    input LPBKRXTXSEREN;
    input LPBKTXRXSEREN;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input QPLL0CLK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RSTCLKENTX;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input RXCOMMADETEN;
    input RXDCCFORCESTART;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input [3:0] RXOSINTCFG;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input [2:0] TXBUFDIFFCTRL;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXELFORCESTART;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTYE3_COMMON (...);
    parameter [15:0] A_SDM1DATA1_0 = 16'b0000000000000000;
    parameter [8:0] A_SDM1DATA1_1 = 9'b000000000;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [9:0] BIAS_CFG_RSVD = 10'b0000000000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0004;
    parameter [15:0] PPF0_CFG = 16'h0FFF;
    parameter [15:0] PPF1_CFG = 16'h0FFF;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h301C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0780;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0780;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0021;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1111111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter integer QPLL0_REFCLK_DIV = 2;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h301C;
    parameter [15:0] QPLL1_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0780;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0780;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0021;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1111111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter integer QPLL1_REFCLK_DIV = 2;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_EN = 1'b1;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer SIM_VERSION = 2;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0_SEL;
    output [1:0] RXRECCLK1_SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input [1:0] SDM1WIDTH;
endmodule

module GTYE4_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_RXTERMINATION = 1'b1;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter [0:0] CFOK_PWRSVE_EN = 1'b1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h2424;
    parameter [15:0] CKCAL1_CFG_0 = 16'b1100000011000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0101000011000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b1100000011000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b1000000011000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h01FA;
    parameter [15:0] CPLL_CFG1 = 16'h24A9;
    parameter [15:0] CPLL_CFG2 = 16'h6807;
    parameter [15:0] CPLL_CFG3 = 16'h0000;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DELAY_ELEC = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h800;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter integer EYESCAN_VP_RANGE = 0;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter integer LPBK_BIAS_CTRL = 4;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter integer LPBK_IND_CTRL0 = 5;
    parameter integer LPBK_IND_CTRL1 = 5;
    parameter integer LPBK_IND_CTRL2 = 5;
    parameter integer LPBK_RG_CTRL = 2;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'b00000;
    parameter [5:0] PCIE3_CLK_COR_FULL_THRSH = 6'b010000;
    parameter [4:0] PCIE3_CLK_COR_MAX_LAT = 5'b01000;
    parameter [4:0] PCIE3_CLK_COR_MIN_LAT = 5'b00100;
    parameter [5:0] PCIE3_CLK_COR_THRSH_TIMER = 6'b001000;
    parameter PCIE_64B_DYN_CLKSW_DIS = "FALSE";
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter PCIE_GEN4_64BIT_INT_EN = "FALSE";
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN4 = 2'h0;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'h0000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0;
    parameter [0:0] RCLK_SIPO_INV_EN = 1'b0;
    parameter [2:0] RTX_BUF_CML_CTRL = 3'b010;
    parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b10000;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0003;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0003;
    parameter [15:0] RXCDR_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h0164;
    parameter [9:0] RXCDR_CFG2_GEN2 = 10'h164;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0034;
    parameter [15:0] RXCDR_CFG2_GEN4 = 16'h0034;
    parameter [15:0] RXCDR_CFG3 = 16'h0024;
    parameter [5:0] RXCDR_CFG3_GEN2 = 6'h24;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0024;
    parameter [15:0] RXCDR_CFG3_GEN4 = 16'h0024;
    parameter [15:0] RXCDR_CFG4 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG5 = 16'hB46B;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h146B;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h0000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0002;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_KH_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG3 = 16'h2000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_UT_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h1000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000110000;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] RXPI_CFG0 = 16'h0102;
    parameter [15:0] RXPI_CFG1 = 16'b0000000001010100;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter [0:0] RXREFCLKDIV2_SEL = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h12B0;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 2;
    parameter integer RX_CM_TRIM = 12;
    parameter [0:0] RX_CTLE_PWR_SAVING = 1'b0;
    parameter [3:0] RX_CTLE_RES_CTRL = 4'b0000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b100;
    parameter integer RX_DFELPM_CFG0 = 10;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b1;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 2;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter integer RX_EN_SUM_RCAL_B = 0;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b10;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] RX_I2V_FILTER_EN = 1'b1;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] RX_PMA_RSV0 = 16'h002F;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter integer RX_SUM_DEGEN_AVTT_OVERITE = 0;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter integer RX_SUM_PWR_SAVING = 0;
    parameter [3:0] RX_SUM_RES_CTRL = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b0011;
    parameter [0:0] RX_SUM_VCM_BIAS_TUNE_EN = 1'b1;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b010;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter [0:0] SAMPLE_CLK_PHASE = 1'b0;
    parameter [0:0] SAS_12G_MODE = 1'b0;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
    parameter [0:0] SRSTMODE = 1'b0;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter integer TXDRV_FREQBAND = 0;
    parameter [15:0] TXFE_CFG0 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG1 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG2 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG3 = 16'b0000000000000000;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h6020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0002;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] TXPI_CFG0 = 16'b0000000100000000;
    parameter [15:0] TXPI_CFG1 = 16'b0000000000000000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_PPM = 1'b0;
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXREFCLKDIV2_SEL = 1'b0;
    parameter integer TXSWBST_BST = 1;
    parameter integer TXSWBST_EN = 0;
    parameter integer TXSWBST_MAG = 6;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [5:0] TX_DEEMPH2 = 6'b000000;
    parameter [5:0] TX_DEEMPH3 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h003F;
    parameter integer TX_PI_BIASSET = 0;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] TX_PMA_RSV0 = 16'h0000;
    parameter [15:0] TX_PMA_RSV1 = 16'h0000;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 3;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [1:0] TX_SW_MEAS = 2'b00;
    parameter [2:0] TX_VREG_CTRL = 3'b000;
    parameter [0:0] TX_VREG_PDB = 1'b0;
    parameter [1:0] TX_VREG_VREFSEL = 2'b00;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USB_BOTH_BURST_IDLE = 1'b0;
    parameter [6:0] USB_BURSTMAX_U3WAKE = 7'b1111111;
    parameter [6:0] USB_BURSTMIN_U3WAKE = 7'b1100011;
    parameter [0:0] USB_CLK_COR_EQ_EN = 1'b0;
    parameter [0:0] USB_EXT_CNTL = 1'b1;
    parameter [9:0] USB_IDLEMAX_POLLING = 10'b1010111011;
    parameter [9:0] USB_IDLEMIN_POLLING = 10'b0100101011;
    parameter [8:0] USB_LFPSPING_BURST = 9'b000000101;
    parameter [8:0] USB_LFPSPOLLING_BURST = 9'b000110001;
    parameter [8:0] USB_LFPSPOLLING_IDLE_MS = 9'b000000100;
    parameter [8:0] USB_LFPSU1EXIT_BURST = 9'b000011101;
    parameter [8:0] USB_LFPSU2LPEXIT_BURST_MS = 9'b001100011;
    parameter [8:0] USB_LFPSU3WAKE_BURST_MS = 9'b111110011;
    parameter [3:0] USB_LFPS_TPERIOD = 4'b0011;
    parameter [0:0] USB_LFPS_TPERIOD_ACCURATE = 1'b1;
    parameter [0:0] USB_MODE = 1'b0;
    parameter [0:0] USB_PCIE_ERR_REP_DIS = 1'b0;
    parameter integer USB_PING_SATA_MAX_INIT = 21;
    parameter integer USB_PING_SATA_MIN_INIT = 12;
    parameter integer USB_POLL_SATA_MAX_BURST = 8;
    parameter integer USB_POLL_SATA_MIN_BURST = 4;
    parameter [0:0] USB_RAW_ELEC = 1'b0;
    parameter [0:0] USB_RXIDLE_P0_CTRL = 1'b1;
    parameter [0:0] USB_TXIDLE_TUNE_ENABLE = 1'b1;
    parameter integer USB_U1_SATA_MAX_WAKE = 7;
    parameter integer USB_U1_SATA_MIN_WAKE = 4;
    parameter integer USB_U2_SAS_MAX_COM = 64;
    parameter integer USB_U2_SAS_MIN_COM = 36;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [0:0] Y_ALL_MODE = 1'b0;
    output BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [15:0] DMONITOROUT;
    output DMONITOROUTCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output GTYTXN;
    output GTYTXP;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [15:0] PINRSRVDAS;
    output POWERPRESENT;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output RXLFPSTRESETDET;
    output RXLFPSU2LPEXITDET;
    output RXLFPSU3WAKEDET;
    output [7:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLFREQLOCK;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input FREQOS;
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTRXRESETSEL;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTTXRESETSEL;
    input GTYRXN;
    input GTYRXP;
    input INCPCTRL;
    input [2:0] LOOPBACK;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input QPLL0CLK;
    input QPLL0FREQLOCK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1FREQLOCK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXAFECFOKEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input [6:0] RXCKCALSTART;
    input RXCOMMADETEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input [3:0] RXDFECFOKFCNUM;
    input RXDFECFOKFEN;
    input RXDFECFOKFPULSE;
    input RXDFECFOKHOLD;
    input RXDFECFOKOVREN;
    input RXDFEKHHOLD;
    input RXDFEKHOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXEQTRAINING;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXTERMINATION;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input [1:0] TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input TXLFPSTRESET;
    input TXLFPSU2LPEXIT;
    input TXLFPSU3WAKE;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input TXMUXDCDEXHOLD;
    input TXMUXDCDORWREN;
    input TXONESZEROS;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTYE4_COMMON (...);
    parameter [0:0] AEN_QPLL0_FBDIV = 1'b1;
    parameter [0:0] AEN_QPLL1_FBDIV = 1'b1;
    parameter [0:0] AEN_SDM0TOGGLE = 1'b0;
    parameter [0:0] AEN_SDM1TOGGLE = 1'b0;
    parameter [0:0] A_SDM0TOGGLE = 1'b0;
    parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000;
    parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000;
    parameter [0:0] A_SDM1TOGGLE = 1'b0;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [15:0] BIAS_CFG_RSVD = 16'h0000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0000;
    parameter [15:0] PPF0_CFG = 16'h0F00;
    parameter [15:0] PPF1_CFG = 16'h0F00;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h391C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0F80;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0002;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1011111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL0_PCI_EN = 1'b0;
    parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL0_REFCLK_DIV = 1;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h691C;
    parameter [15:0] QPLL1_CFG1 = 16'h0020;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0F80;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0002;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1011111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL1_PCI_EN = 1'b0;
    parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL1_REFCLK_DIV = 1;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_ENB = 1'b0;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [15:0] UB_CFG0 = 16'h0000;
    parameter [15:0] UB_CFG1 = 16'h0000;
    parameter [15:0] UB_CFG2 = 16'h0000;
    parameter [15:0] UB_CFG3 = 16'h0000;
    parameter [15:0] UB_CFG4 = 16'h0000;
    parameter [15:0] UB_CFG5 = 16'h0400;
    parameter [15:0] UB_CFG6 = 16'h0000;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0SEL;
    output [1:0] RXRECCLK1SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    output [15:0] UBDADDR;
    output UBDEN;
    output [15:0] UBDI;
    output UBDWE;
    output UBMDMTDO;
    output UBRSVDOUT;
    output UBTXUART;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [15:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [2:0] PCIERATEQPLL0;
    input [2:0] PCIERATEQPLL1;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input [7:0] QPLL0FBDIV;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input [7:0] QPLL1FBDIV;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input SDM0TOGGLE;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input SDM1TOGGLE;
    input [1:0] SDM1WIDTH;
    input UBCFGSTREAMEN;
    input [15:0] UBDO;
    input UBDRDY;
    input UBENABLE;
    input [1:0] UBGPI;
    input [1:0] UBINTR;
    input UBIOLMBRST;
    input UBMBRST;
    input UBMDMCAPTURE;
    input UBMDMDBGRST;
    input UBMDMDBGUPDATE;
    input [3:0] UBMDMREGEN;
    input UBMDMSHIFT;
    input UBMDMSYSRST;
    input UBMDMTCK;
    input UBMDMTDI;
endmodule

module IBUFDS_GTE3 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [1:0] REFCLK_HROW_CK_SEL = 2'b00;
    parameter [1:0] REFCLK_ICNTL_RX = 2'b00;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_GTE4 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [1:0] REFCLK_HROW_CK_SEL = 2'b00;
    parameter [1:0] REFCLK_ICNTL_RX = 2'b00;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module OBUFDS_GTE3 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTE3_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
    input [1:0] RXRECCLK_SEL;
endmodule

module OBUFDS_GTE4 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTE4_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
    input [1:0] RXRECCLK_SEL;
endmodule

module PCIE_A1 (...);
    parameter [31:0] BAR0 = 32'h00000000;
    parameter [31:0] BAR1 = 32'h00000000;
    parameter [31:0] BAR2 = 32'h00000000;
    parameter [31:0] BAR3 = 32'h00000000;
    parameter [31:0] BAR4 = 32'h00000000;
    parameter [31:0] BAR5 = 32'h00000000;
    parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
    parameter [23:0] CLASS_CODE = 24'h000000;
    parameter integer DEV_CAP_ENDPOINT_L0S_LATENCY = 7;
    parameter integer DEV_CAP_ENDPOINT_L1_LATENCY = 7;
    parameter DEV_CAP_EXT_TAG_SUPPORTED = "FALSE";
    parameter integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
    parameter integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
    parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
    parameter DISABLE_BAR_FILTERING = "FALSE";
    parameter DISABLE_ID_CHECK = "FALSE";
    parameter DISABLE_SCRAMBLING = "FALSE";
    parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
    parameter [21:0] EXPANSION_ROM = 22'h000000;
    parameter FAST_TRAIN = "FALSE";
    parameter integer GTP_SEL = 0;
    parameter integer LINK_CAP_ASPM_SUPPORT = 1;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY = 7;
    parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "FALSE";
    parameter [14:0] LL_ACK_TIMEOUT = 15'h0204;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter [14:0] LL_REPLAY_TIMEOUT = 15'h060D;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer MSI_CAP_MULTIMSGCAP = 0;
    parameter integer MSI_CAP_MULTIMSG_EXTENSION = 0;
    parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h1;
    parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
    parameter [4:0] PCIE_CAP_INT_MSG_NUM = 5'b00000;
    parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
    parameter [11:0] PCIE_GENERIC = 12'h000;
    parameter PLM_AUTO_CONFIG = "FALSE";
    parameter integer PM_CAP_AUXCURRENT = 0;
    parameter PM_CAP_D1SUPPORT = "TRUE";
    parameter PM_CAP_D2SUPPORT = "TRUE";
    parameter PM_CAP_DSI = "FALSE";
    parameter [4:0] PM_CAP_PMESUPPORT = 5'b01111;
    parameter PM_CAP_PME_CLOCK = "FALSE";
    parameter integer PM_CAP_VERSION = 3;
    parameter [7:0] PM_DATA0 = 8'h1E;
    parameter [7:0] PM_DATA1 = 8'h1E;
    parameter [7:0] PM_DATA2 = 8'h1E;
    parameter [7:0] PM_DATA3 = 8'h1E;
    parameter [7:0] PM_DATA4 = 8'h1E;
    parameter [7:0] PM_DATA5 = 8'h1E;
    parameter [7:0] PM_DATA6 = 8'h1E;
    parameter [7:0] PM_DATA7 = 8'h1E;
    parameter [1:0] PM_DATA_SCALE0 = 2'b01;
    parameter [1:0] PM_DATA_SCALE1 = 2'b01;
    parameter [1:0] PM_DATA_SCALE2 = 2'b01;
    parameter [1:0] PM_DATA_SCALE3 = 2'b01;
    parameter [1:0] PM_DATA_SCALE4 = 2'b01;
    parameter [1:0] PM_DATA_SCALE5 = 2'b01;
    parameter [1:0] PM_DATA_SCALE6 = 2'b01;
    parameter [1:0] PM_DATA_SCALE7 = 2'b01;
    parameter SIM_VERSION = "1.0";
    parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
    parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
    parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
    parameter integer TL_RX_RAM_RADDR_LATENCY = 1;
    parameter integer TL_RX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_RX_RAM_WRITE_LATENCY = 0;
    parameter TL_TFC_DISABLE = "FALSE";
    parameter TL_TX_CHECKS_DISABLE = "FALSE";
    parameter integer TL_TX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_TX_RAM_RDATA_LATENCY = 2;
    parameter USR_CFG = "FALSE";
    parameter USR_EXT_CFG = "FALSE";
    parameter VC0_CPL_INFINITE = "TRUE";
    parameter [11:0] VC0_RX_RAM_LIMIT = 12'h01E;
    parameter integer VC0_TOTAL_CREDITS_CD = 104;
    parameter integer VC0_TOTAL_CREDITS_CH = 36;
    parameter integer VC0_TOTAL_CREDITS_NPH = 8;
    parameter integer VC0_TOTAL_CREDITS_PD = 288;
    parameter integer VC0_TOTAL_CREDITS_PH = 32;
    parameter integer VC0_TX_LASTPACKET = 31;
    output CFGCOMMANDBUSMASTERENABLE;
    output CFGCOMMANDINTERRUPTDISABLE;
    output CFGCOMMANDIOENABLE;
    output CFGCOMMANDMEMENABLE;
    output CFGCOMMANDSERREN;
    output CFGDEVCONTROLAUXPOWEREN;
    output CFGDEVCONTROLCORRERRREPORTINGEN;
    output CFGDEVCONTROLENABLERO;
    output CFGDEVCONTROLEXTTAGEN;
    output CFGDEVCONTROLFATALERRREPORTINGEN;
    output CFGDEVCONTROLNONFATALREPORTINGEN;
    output CFGDEVCONTROLNOSNOOPEN;
    output CFGDEVCONTROLPHANTOMEN;
    output CFGDEVCONTROLURERRREPORTINGEN;
    output CFGDEVSTATUSCORRERRDETECTED;
    output CFGDEVSTATUSFATALERRDETECTED;
    output CFGDEVSTATUSNONFATALERRDETECTED;
    output CFGDEVSTATUSURDETECTED;
    output CFGERRCPLRDYN;
    output CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTRDYN;
    output CFGLINKCONTOLRCB;
    output CFGLINKCONTROLCOMMONCLOCK;
    output CFGLINKCONTROLEXTENDEDSYNC;
    output CFGRDWRDONEN;
    output CFGTOTURNOFFN;
    output DBGBADDLLPSTATUS;
    output DBGBADTLPLCRC;
    output DBGBADTLPSEQNUM;
    output DBGBADTLPSTATUS;
    output DBGDLPROTOCOLSTATUS;
    output DBGFCPROTOCOLERRSTATUS;
    output DBGMLFRMDLENGTH;
    output DBGMLFRMDMPS;
    output DBGMLFRMDTCVC;
    output DBGMLFRMDTLPSTATUS;
    output DBGMLFRMDUNRECTYPE;
    output DBGPOISTLPSTATUS;
    output DBGRCVROVERFLOWSTATUS;
    output DBGREGDETECTEDCORRECTABLE;
    output DBGREGDETECTEDFATAL;
    output DBGREGDETECTEDNONFATAL;
    output DBGREGDETECTEDUNSUPPORTED;
    output DBGRPLYROLLOVERSTATUS;
    output DBGRPLYTIMEOUTSTATUS;
    output DBGURNOBARHIT;
    output DBGURPOISCFGWR;
    output DBGURSTATUS;
    output DBGURUNSUPMSG;
    output MIMRXREN;
    output MIMRXWEN;
    output MIMTXREN;
    output MIMTXWEN;
    output PIPEGTTXELECIDLEA;
    output PIPEGTTXELECIDLEB;
    output PIPERXPOLARITYA;
    output PIPERXPOLARITYB;
    output PIPERXRESETA;
    output PIPERXRESETB;
    output PIPETXRCVRDETA;
    output PIPETXRCVRDETB;
    output RECEIVEDHOTRESET;
    output TRNLNKUPN;
    output TRNREOFN;
    output TRNRERRFWDN;
    output TRNRSOFN;
    output TRNRSRCDSCN;
    output TRNRSRCRDYN;
    output TRNTCFGREQN;
    output TRNTDSTRDYN;
    output TRNTERRDROPN;
    output USERRSTN;
    output [11:0] MIMRXRADDR;
    output [11:0] MIMRXWADDR;
    output [11:0] MIMTXRADDR;
    output [11:0] MIMTXWADDR;
    output [11:0] TRNFCCPLD;
    output [11:0] TRNFCNPD;
    output [11:0] TRNFCPD;
    output [15:0] PIPETXDATAA;
    output [15:0] PIPETXDATAB;
    output [1:0] CFGLINKCONTROLASPMCONTROL;
    output [1:0] PIPEGTPOWERDOWNA;
    output [1:0] PIPEGTPOWERDOWNB;
    output [1:0] PIPETXCHARDISPMODEA;
    output [1:0] PIPETXCHARDISPMODEB;
    output [1:0] PIPETXCHARDISPVALA;
    output [1:0] PIPETXCHARDISPVALB;
    output [1:0] PIPETXCHARISKA;
    output [1:0] PIPETXCHARISKB;
    output [2:0] CFGDEVCONTROLMAXPAYLOAD;
    output [2:0] CFGDEVCONTROLMAXREADREQ;
    output [2:0] CFGFUNCTIONNUMBER;
    output [2:0] CFGINTERRUPTMMENABLE;
    output [2:0] CFGPCIELINKSTATEN;
    output [31:0] CFGDO;
    output [31:0] TRNRD;
    output [34:0] MIMRXWDATA;
    output [35:0] MIMTXWDATA;
    output [4:0] CFGDEVICENUMBER;
    output [4:0] CFGLTSSMSTATE;
    output [5:0] TRNTBUFAV;
    output [6:0] TRNRBARHITN;
    output [7:0] CFGBUSNUMBER;
    output [7:0] CFGINTERRUPTDO;
    output [7:0] TRNFCCPLH;
    output [7:0] TRNFCNPH;
    output [7:0] TRNFCPH;
    input CFGERRCORN;
    input CFGERRCPLABORTN;
    input CFGERRCPLTIMEOUTN;
    input CFGERRECRCN;
    input CFGERRLOCKEDN;
    input CFGERRPOSTEDN;
    input CFGERRURN;
    input CFGINTERRUPTASSERTN;
    input CFGINTERRUPTN;
    input CFGPMWAKEN;
    input CFGRDENN;
    input CFGTRNPENDINGN;
    input CFGTURNOFFOKN;
    input CLOCKLOCKED;
    input MGTCLK;
    input PIPEGTRESETDONEA;
    input PIPEGTRESETDONEB;
    input PIPEPHYSTATUSA;
    input PIPEPHYSTATUSB;
    input PIPERXENTERELECIDLEA;
    input PIPERXENTERELECIDLEB;
    input SYSRESETN;
    input TRNRDSTRDYN;
    input TRNRNPOKN;
    input TRNTCFGGNTN;
    input TRNTEOFN;
    input TRNTERRFWDN;
    input TRNTSOFN;
    input TRNTSRCDSCN;
    input TRNTSRCRDYN;
    input TRNTSTRN;
    input USERCLK;
    input [15:0] CFGDEVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENID;
    input [15:0] CFGVENID;
    input [15:0] PIPERXDATAA;
    input [15:0] PIPERXDATAB;
    input [1:0] PIPERXCHARISKA;
    input [1:0] PIPERXCHARISKB;
    input [2:0] PIPERXSTATUSA;
    input [2:0] PIPERXSTATUSB;
    input [2:0] TRNFCSEL;
    input [31:0] TRNTD;
    input [34:0] MIMRXRDATA;
    input [35:0] MIMTXRDATA;
    input [47:0] CFGERRTLPCPLHEADER;
    input [63:0] CFGDSN;
    input [7:0] CFGINTERRUPTDI;
    input [7:0] CFGREVID;
    input [9:0] CFGDWADDR;
endmodule

module PCIE_EP (...);
    parameter BAR0EXIST = "TRUE";
    parameter BAR0PREFETCHABLE = "TRUE";
    parameter BAR1EXIST = "FALSE";
    parameter BAR1PREFETCHABLE = "FALSE";
    parameter BAR2EXIST = "FALSE";
    parameter BAR2PREFETCHABLE = "FALSE";
    parameter BAR3EXIST = "FALSE";
    parameter BAR3PREFETCHABLE = "FALSE";
    parameter BAR4EXIST = "FALSE";
    parameter BAR4PREFETCHABLE = "FALSE";
    parameter BAR5EXIST = "FALSE";
    parameter BAR5PREFETCHABLE = "FALSE";
    parameter CLKDIVIDED = "FALSE";
    parameter INFINITECOMPLETIONS = "TRUE";
    parameter LINKSTATUSSLOTCLOCKCONFIG = "FALSE";
    parameter PBCAPABILITYSYSTEMALLOCATED = "FALSE";
    parameter PMCAPABILITYD1SUPPORT = "FALSE";
    parameter PMCAPABILITYD2SUPPORT = "FALSE";
    parameter PMCAPABILITYDSI = "TRUE";
    parameter RESETMODE = "FALSE";
    parameter [10:0] VC0TOTALCREDITSCD = 11'h0;
    parameter [10:0] VC0TOTALCREDITSPD = 11'h34;
    parameter [10:0] VC1TOTALCREDITSCD = 11'h0;
    parameter [10:0] VC1TOTALCREDITSPD = 11'h0;
    parameter [11:0] AERBASEPTR = 12'h110;
    parameter [11:0] AERCAPABILITYNEXTPTR = 12'h138;
    parameter [11:0] DSNBASEPTR = 12'h148;
    parameter [11:0] DSNCAPABILITYNEXTPTR = 12'h154;
    parameter [11:0] MSIBASEPTR = 12'h48;
    parameter [11:0] PBBASEPTR = 12'h138;
    parameter [11:0] PBCAPABILITYNEXTPTR = 12'h148;
    parameter [11:0] PMBASEPTR = 12'h40;
    parameter [11:0] RETRYRAMSIZE = 12'h9;
    parameter [11:0] VCBASEPTR = 12'h154;
    parameter [11:0] VCCAPABILITYNEXTPTR = 12'h0;
    parameter [12:0] VC0RXFIFOBASEC = 13'h98;
    parameter [12:0] VC0RXFIFOBASENP = 13'h80;
    parameter [12:0] VC0RXFIFOBASEP = 13'h0;
    parameter [12:0] VC0RXFIFOLIMITC = 13'h117;
    parameter [12:0] VC0RXFIFOLIMITNP = 13'h97;
    parameter [12:0] VC0RXFIFOLIMITP = 13'h7f;
    parameter [12:0] VC0TXFIFOBASEC = 13'h98;
    parameter [12:0] VC0TXFIFOBASENP = 13'h80;
    parameter [12:0] VC0TXFIFOBASEP = 13'h0;
    parameter [12:0] VC0TXFIFOLIMITC = 13'h117;
    parameter [12:0] VC0TXFIFOLIMITNP = 13'h97;
    parameter [12:0] VC0TXFIFOLIMITP = 13'h7f;
    parameter [12:0] VC1RXFIFOBASEC = 13'h118;
    parameter [12:0] VC1RXFIFOBASENP = 13'h118;
    parameter [12:0] VC1RXFIFOBASEP = 13'h118;
    parameter [12:0] VC1RXFIFOLIMITC = 13'h118;
    parameter [12:0] VC1RXFIFOLIMITNP = 13'h118;
    parameter [12:0] VC1RXFIFOLIMITP = 13'h118;
    parameter [12:0] VC1TXFIFOBASEC = 13'h118;
    parameter [12:0] VC1TXFIFOBASENP = 13'h118;
    parameter [12:0] VC1TXFIFOBASEP = 13'h118;
    parameter [12:0] VC1TXFIFOLIMITC = 13'h118;
    parameter [12:0] VC1TXFIFOLIMITNP = 13'h118;
    parameter [12:0] VC1TXFIFOLIMITP = 13'h118;
    parameter [15:0] DEVICEID = 16'h5050;
    parameter [15:0] SUBSYSTEMID = 16'h5050;
    parameter [15:0] SUBSYSTEMVENDORID = 16'h10EE;
    parameter [15:0] VENDORID = 16'h10EE;
    parameter [1:0] LINKCAPABILITYASPMSUPPORT = 2'h1;
    parameter [1:0] PBCAPABILITYDW0DATASCALE = 2'h0;
    parameter [1:0] PBCAPABILITYDW0PMSTATE = 2'h0;
    parameter [1:0] PBCAPABILITYDW1DATASCALE = 2'h0;
    parameter [1:0] PBCAPABILITYDW1PMSTATE = 2'h0;
    parameter [1:0] PBCAPABILITYDW2DATASCALE = 2'h0;
    parameter [1:0] PBCAPABILITYDW2PMSTATE = 2'h0;
    parameter [1:0] PBCAPABILITYDW3DATASCALE = 2'h0;
    parameter [1:0] PBCAPABILITYDW3PMSTATE = 2'h0;
    parameter [23:0] CLASSCODE = 24'h058000;
    parameter [2:0] DEVICECAPABILITYENDPOINTL0SLATENCY = 3'h0;
    parameter [2:0] DEVICECAPABILITYENDPOINTL1LATENCY = 3'h0;
    parameter [2:0] MSICAPABILITYMULTIMSGCAP = 3'h0;
    parameter [2:0] PBCAPABILITYDW0PMSUBSTATE = 3'h0;
    parameter [2:0] PBCAPABILITYDW0POWERRAIL = 3'h0;
    parameter [2:0] PBCAPABILITYDW0TYPE = 3'h0;
    parameter [2:0] PBCAPABILITYDW1PMSUBSTATE = 3'h0;
    parameter [2:0] PBCAPABILITYDW1POWERRAIL = 3'h0;
    parameter [2:0] PBCAPABILITYDW1TYPE = 3'h0;
    parameter [2:0] PBCAPABILITYDW2PMSUBSTATE = 3'h0;
    parameter [2:0] PBCAPABILITYDW2POWERRAIL = 3'h0;
    parameter [2:0] PBCAPABILITYDW2TYPE = 3'h0;
    parameter [2:0] PBCAPABILITYDW3PMSUBSTATE = 3'h0;
    parameter [2:0] PBCAPABILITYDW3POWERRAIL = 3'h0;
    parameter [2:0] PBCAPABILITYDW3TYPE = 3'h0;
    parameter [2:0] PMCAPABILITYAUXCURRENT = 3'h0;
    parameter [2:0] PORTVCCAPABILITYEXTENDEDVCCOUNT = 3'h0;
    parameter [31:0] CARDBUSCISPOINTER = 32'h0;
    parameter [3:0] XPDEVICEPORTTYPE = 4'h0;
    parameter [4:0] PMCAPABILITYPMESUPPORT = 5'h0;
    parameter [5:0] BAR0MASKWIDTH = 6'h14;
    parameter [5:0] BAR1MASKWIDTH = 6'h0;
    parameter [5:0] BAR2MASKWIDTH = 6'h0;
    parameter [5:0] BAR3MASKWIDTH = 6'h0;
    parameter [5:0] BAR4MASKWIDTH = 6'h0;
    parameter [5:0] BAR5MASKWIDTH = 6'h0;
    parameter [5:0] LINKCAPABILITYMAXLINKWIDTH = 6'h01;
    parameter [63:0] DEVICESERIALNUMBER = 64'hE000000001000A35;
    parameter [6:0] VC0TOTALCREDITSCH = 7'h0;
    parameter [6:0] VC0TOTALCREDITSNPH = 7'h08;
    parameter [6:0] VC0TOTALCREDITSPH = 7'h08;
    parameter [6:0] VC1TOTALCREDITSCH = 7'h0;
    parameter [6:0] VC1TOTALCREDITSNPH = 7'h0;
    parameter [6:0] VC1TOTALCREDITSPH = 7'h0;
    parameter [7:0] ACTIVELANESIN = 8'h1;
    parameter [7:0] CAPABILITIESPOINTER = 8'h40;
    parameter [7:0] INTERRUPTPIN = 8'h0;
    parameter [7:0] MSICAPABILITYNEXTPTR = 8'h60;
    parameter [7:0] PBCAPABILITYDW0BASEPOWER = 8'h0;
    parameter [7:0] PBCAPABILITYDW1BASEPOWER = 8'h0;
    parameter [7:0] PBCAPABILITYDW2BASEPOWER = 8'h0;
    parameter [7:0] PBCAPABILITYDW3BASEPOWER = 8'h0;
    parameter [7:0] PCIECAPABILITYNEXTPTR = 8'h0;
    parameter [7:0] PMCAPABILITYNEXTPTR = 8'h60;
    parameter [7:0] PMDATA0 = 8'h0;
    parameter [7:0] PMDATA1 = 8'h0;
    parameter [7:0] PMDATA2 = 8'h0;
    parameter [7:0] PMDATA3 = 8'h0;
    parameter [7:0] PMDATA4 = 8'h0;
    parameter [7:0] PMDATA5 = 8'h0;
    parameter [7:0] PMDATA6 = 8'h0;
    parameter [7:0] PMDATA7 = 8'h0;
    parameter [7:0] PORTVCCAPABILITYVCARBCAP = 8'h0;
    parameter [7:0] PORTVCCAPABILITYVCARBTABLEOFFSET = 8'h0;
    parameter [7:0] REVISIONID = 8'h0;
    parameter [7:0] XPBASEPTR = 8'h60;
    parameter BAR0ADDRWIDTH = 0;
    parameter BAR0IOMEMN = 0;
    parameter BAR1ADDRWIDTH = 0;
    parameter BAR1IOMEMN = 0;
    parameter BAR2ADDRWIDTH = 0;
    parameter BAR2IOMEMN = 0;
    parameter BAR3ADDRWIDTH = 0;
    parameter BAR3IOMEMN = 0;
    parameter BAR4ADDRWIDTH = 0;
    parameter BAR4IOMEMN = 0;
    parameter BAR5IOMEMN = 0;
    parameter L0SEXITLATENCY = 7;
    parameter L0SEXITLATENCYCOMCLK = 7;
    parameter L1EXITLATENCY = 7;
    parameter L1EXITLATENCYCOMCLK = 7;
    parameter LOWPRIORITYVCCOUNT = 0;
    parameter PMDATASCALE0 = 0;
    parameter PMDATASCALE1 = 0;
    parameter PMDATASCALE2 = 0;
    parameter PMDATASCALE3 = 0;
    parameter PMDATASCALE4 = 0;
    parameter PMDATASCALE5 = 0;
    parameter PMDATASCALE6 = 0;
    parameter PMDATASCALE7 = 0;
    parameter RETRYRAMREADLATENCY = 3;
    parameter RETRYRAMWRITELATENCY = 1;
    parameter TLRAMREADLATENCY = 3;
    parameter TLRAMWRITELATENCY = 1;
    parameter TXTSNFTS = 255;
    parameter TXTSNFTSCOMCLK = 255;
    parameter XPMAXPAYLOAD = 0;
    output BUSMASTERENABLE;
    output CRMDOHOTRESETN;
    output CRMPWRSOFTRESETN;
    output DLLTXPMDLLPOUTSTANDING;
    output INTERRUPTDISABLE;
    output IOSPACEENABLE;
    output L0CFGLOOPBACKACK;
    output L0DLLRXACKOUTSTANDING;
    output L0DLLTXNONFCOUTSTANDING;
    output L0DLLTXOUTSTANDING;
    output L0FIRSTCFGWRITEOCCURRED;
    output L0MACENTEREDL0;
    output L0MACLINKTRAINING;
    output L0MACLINKUP;
    output L0MACNEWSTATEACK;
    output L0MACRXL0SSTATE;
    output L0MSIENABLE0;
    output L0PMEACK;
    output L0PMEEN;
    output L0PMEREQOUT;
    output L0PWRL1STATE;
    output L0PWRL23READYSTATE;
    output L0PWRTURNOFFREQ;
    output L0PWRTXL0SSTATE;
    output L0RXDLLPM;
    output L0STATSCFGOTHERRECEIVED;
    output L0STATSCFGOTHERTRANSMITTED;
    output L0STATSCFGRECEIVED;
    output L0STATSCFGTRANSMITTED;
    output L0STATSDLLPRECEIVED;
    output L0STATSDLLPTRANSMITTED;
    output L0STATSOSRECEIVED;
    output L0STATSOSTRANSMITTED;
    output L0STATSTLPRECEIVED;
    output L0STATSTLPTRANSMITTED;
    output L0UNLOCKRECEIVED;
    output LLKRXEOFN;
    output LLKRXEOPN;
    output LLKRXSOFN;
    output LLKRXSOPN;
    output LLKRXSRCLASTREQN;
    output LLKRXSRCRDYN;
    output LLKTXCONFIGREADYN;
    output LLKTXDSTRDYN;
    output MEMSPACEENABLE;
    output MIMDLLBREN;
    output MIMDLLBWEN;
    output MIMRXBREN;
    output MIMRXBWEN;
    output MIMTXBREN;
    output MIMTXBWEN;
    output PARITYERRORRESPONSE;
    output PIPEDESKEWLANESL0;
    output PIPEDESKEWLANESL1;
    output PIPEDESKEWLANESL2;
    output PIPEDESKEWLANESL3;
    output PIPEDESKEWLANESL4;
    output PIPEDESKEWLANESL5;
    output PIPEDESKEWLANESL6;
    output PIPEDESKEWLANESL7;
    output PIPERESETL0;
    output PIPERESETL1;
    output PIPERESETL2;
    output PIPERESETL3;
    output PIPERESETL4;
    output PIPERESETL5;
    output PIPERESETL6;
    output PIPERESETL7;
    output PIPERXPOLARITYL0;
    output PIPERXPOLARITYL1;
    output PIPERXPOLARITYL2;
    output PIPERXPOLARITYL3;
    output PIPERXPOLARITYL4;
    output PIPERXPOLARITYL5;
    output PIPERXPOLARITYL6;
    output PIPERXPOLARITYL7;
    output PIPETXCOMPLIANCEL0;
    output PIPETXCOMPLIANCEL1;
    output PIPETXCOMPLIANCEL2;
    output PIPETXCOMPLIANCEL3;
    output PIPETXCOMPLIANCEL4;
    output PIPETXCOMPLIANCEL5;
    output PIPETXCOMPLIANCEL6;
    output PIPETXCOMPLIANCEL7;
    output PIPETXDATAKL0;
    output PIPETXDATAKL1;
    output PIPETXDATAKL2;
    output PIPETXDATAKL3;
    output PIPETXDATAKL4;
    output PIPETXDATAKL5;
    output PIPETXDATAKL6;
    output PIPETXDATAKL7;
    output PIPETXDETECTRXLOOPBACKL0;
    output PIPETXDETECTRXLOOPBACKL1;
    output PIPETXDETECTRXLOOPBACKL2;
    output PIPETXDETECTRXLOOPBACKL3;
    output PIPETXDETECTRXLOOPBACKL4;
    output PIPETXDETECTRXLOOPBACKL5;
    output PIPETXDETECTRXLOOPBACKL6;
    output PIPETXDETECTRXLOOPBACKL7;
    output PIPETXELECIDLEL0;
    output PIPETXELECIDLEL1;
    output PIPETXELECIDLEL2;
    output PIPETXELECIDLEL3;
    output PIPETXELECIDLEL4;
    output PIPETXELECIDLEL5;
    output PIPETXELECIDLEL6;
    output PIPETXELECIDLEL7;
    output SERRENABLE;
    output URREPORTINGENABLE;
    output [11:0] MGMTSTATSCREDIT;
    output [11:0] MIMDLLBRADD;
    output [11:0] MIMDLLBWADD;
    output [12:0] L0COMPLETERID;
    output [12:0] MIMRXBRADD;
    output [12:0] MIMRXBWADD;
    output [12:0] MIMTXBRADD;
    output [12:0] MIMTXBWADD;
    output [15:0] LLKRXPREFERREDTYPE;
    output [16:0] MGMTPSO;
    output [1:0] L0PWRSTATE0;
    output [1:0] L0RXMACLINKERROR;
    output [1:0] LLKRXVALIDN;
    output [1:0] PIPEPOWERDOWNL0;
    output [1:0] PIPEPOWERDOWNL1;
    output [1:0] PIPEPOWERDOWNL2;
    output [1:0] PIPEPOWERDOWNL3;
    output [1:0] PIPEPOWERDOWNL4;
    output [1:0] PIPEPOWERDOWNL5;
    output [1:0] PIPEPOWERDOWNL6;
    output [1:0] PIPEPOWERDOWNL7;
    output [2:0] L0MULTIMSGEN0;
    output [2:0] L0RXDLLPMTYPE;
    output [2:0] MAXPAYLOADSIZE;
    output [2:0] MAXREADREQUESTSIZE;
    output [31:0] MGMTRDATA;
    output [3:0] L0LTSSMSTATE;
    output [3:0] L0MACNEGOTIATEDLINKWIDTH;
    output [63:0] LLKRXDATA;
    output [63:0] MIMDLLBWDATA;
    output [63:0] MIMRXBWDATA;
    output [63:0] MIMTXBWDATA;
    output [6:0] L0DLLERRORVECTOR;
    output [7:0] L0DLLVCSTATUS;
    output [7:0] L0DLUPDOWN;
    output [7:0] LLKRXCHCOMPLETIONAVAILABLEN;
    output [7:0] LLKRXCHNONPOSTEDAVAILABLEN;
    output [7:0] LLKRXCHPOSTEDAVAILABLEN;
    output [7:0] LLKTCSTATUS;
    output [7:0] LLKTXCHCOMPLETIONREADYN;
    output [7:0] LLKTXCHNONPOSTEDREADYN;
    output [7:0] LLKTXCHPOSTEDREADYN;
    output [7:0] PIPETXDATAL0;
    output [7:0] PIPETXDATAL1;
    output [7:0] PIPETXDATAL2;
    output [7:0] PIPETXDATAL3;
    output [7:0] PIPETXDATAL4;
    output [7:0] PIPETXDATAL5;
    output [7:0] PIPETXDATAL6;
    output [7:0] PIPETXDATAL7;
    output [9:0] LLKTXCHANSPACE;
    input AUXPOWER;
    input COMPLIANCEAVOID;
    input CRMCORECLK;
    input CRMCORECLKDLO;
    input CRMCORECLKRXO;
    input CRMCORECLKTXO;
    input CRMLINKRSTN;
    input CRMMACRSTN;
    input CRMMGMTRSTN;
    input CRMNVRSTN;
    input CRMURSTN;
    input CRMUSERCFGRSTN;
    input CRMUSERCLK;
    input CRMUSERCLKRXO;
    input CRMUSERCLKTXO;
    input L0CFGDISABLESCRAMBLE;
    input L0CFGLOOPBACKMASTER;
    input L0LEGACYINTFUNCT0;
    input L0PMEREQIN;
    input L0SETCOMPLETERABORTERROR;
    input L0SETCOMPLETIONTIMEOUTCORRERROR;
    input L0SETCOMPLETIONTIMEOUTUNCORRERROR;
    input L0SETDETECTEDCORRERROR;
    input L0SETDETECTEDFATALERROR;
    input L0SETDETECTEDNONFATALERROR;
    input L0SETUNEXPECTEDCOMPLETIONCORRERROR;
    input L0SETUNEXPECTEDCOMPLETIONUNCORRERROR;
    input L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR;
    input L0SETUNSUPPORTEDREQUESTOTHERERROR;
    input L0SETUSERDETECTEDPARITYERROR;
    input L0SETUSERMASTERDATAPARITY;
    input L0SETUSERRECEIVEDMASTERABORT;
    input L0SETUSERRECEIVEDTARGETABORT;
    input L0SETUSERSIGNALLEDTARGETABORT;
    input L0SETUSERSYSTEMERROR;
    input L0TRANSACTIONSPENDING;
    input LLKRXDSTCONTREQN;
    input LLKRXDSTREQN;
    input LLKTXEOFN;
    input LLKTXEOPN;
    input LLKTXSOFN;
    input LLKTXSOPN;
    input LLKTXSRCDSCN;
    input LLKTXSRCRDYN;
    input MGMTRDEN;
    input MGMTWREN;
    input PIPEPHYSTATUSL0;
    input PIPEPHYSTATUSL1;
    input PIPEPHYSTATUSL2;
    input PIPEPHYSTATUSL3;
    input PIPEPHYSTATUSL4;
    input PIPEPHYSTATUSL5;
    input PIPEPHYSTATUSL6;
    input PIPEPHYSTATUSL7;
    input PIPERXCHANISALIGNEDL0;
    input PIPERXCHANISALIGNEDL1;
    input PIPERXCHANISALIGNEDL2;
    input PIPERXCHANISALIGNEDL3;
    input PIPERXCHANISALIGNEDL4;
    input PIPERXCHANISALIGNEDL5;
    input PIPERXCHANISALIGNEDL6;
    input PIPERXCHANISALIGNEDL7;
    input PIPERXDATAKL0;
    input PIPERXDATAKL1;
    input PIPERXDATAKL2;
    input PIPERXDATAKL3;
    input PIPERXDATAKL4;
    input PIPERXDATAKL5;
    input PIPERXDATAKL6;
    input PIPERXDATAKL7;
    input PIPERXELECIDLEL0;
    input PIPERXELECIDLEL1;
    input PIPERXELECIDLEL2;
    input PIPERXELECIDLEL3;
    input PIPERXELECIDLEL4;
    input PIPERXELECIDLEL5;
    input PIPERXELECIDLEL6;
    input PIPERXELECIDLEL7;
    input PIPERXVALIDL0;
    input PIPERXVALIDL1;
    input PIPERXVALIDL2;
    input PIPERXVALIDL3;
    input PIPERXVALIDL4;
    input PIPERXVALIDL5;
    input PIPERXVALIDL6;
    input PIPERXVALIDL7;
    input [10:0] MGMTADDR;
    input [127:0] L0PACKETHEADERFROMUSER;
    input [1:0] LLKRXCHFIFO;
    input [1:0] LLKTXCHFIFO;
    input [1:0] LLKTXENABLEN;
    input [2:0] LLKRXCHTC;
    input [2:0] LLKTXCHTC;
    input [2:0] PIPERXSTATUSL0;
    input [2:0] PIPERXSTATUSL1;
    input [2:0] PIPERXSTATUSL2;
    input [2:0] PIPERXSTATUSL3;
    input [2:0] PIPERXSTATUSL4;
    input [2:0] PIPERXSTATUSL5;
    input [2:0] PIPERXSTATUSL6;
    input [2:0] PIPERXSTATUSL7;
    input [31:0] MGMTWDATA;
    input [3:0] L0MSIREQUEST0;
    input [3:0] MGMTBWREN;
    input [63:0] LLKTXDATA;
    input [63:0] MIMDLLBRDATA;
    input [63:0] MIMRXBRDATA;
    input [63:0] MIMTXBRDATA;
    input [6:0] MGMTSTATSCREDITSEL;
    input [7:0] PIPERXDATAL0;
    input [7:0] PIPERXDATAL1;
    input [7:0] PIPERXDATAL2;
    input [7:0] PIPERXDATAL3;
    input [7:0] PIPERXDATAL4;
    input [7:0] PIPERXDATAL5;
    input [7:0] PIPERXDATAL6;
    input [7:0] PIPERXDATAL7;
endmodule

module PCIE_2_0 (...);
    parameter [11:0] AER_BASE_PTR = 12'h128;
    parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [15:0] AER_CAP_ID = 16'h0001;
    parameter [4:0] AER_CAP_INT_MSG_NUM_MSI = 5'h0A;
    parameter [4:0] AER_CAP_INT_MSG_NUM_MSIX = 5'h15;
    parameter [11:0] AER_CAP_NEXTPTR = 12'h160;
    parameter AER_CAP_ON = "FALSE";
    parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
    parameter [3:0] AER_CAP_VERSION = 4'h1;
    parameter ALLOW_X8_GEN2 = "FALSE";
    parameter [31:0] BAR0 = 32'hFFFFFF00;
    parameter [31:0] BAR1 = 32'hFFFF0000;
    parameter [31:0] BAR2 = 32'hFFFF000C;
    parameter [31:0] BAR3 = 32'hFFFFFFFF;
    parameter [31:0] BAR4 = 32'h00000000;
    parameter [31:0] BAR5 = 32'h00000000;
    parameter [7:0] CAPABILITIES_PTR = 8'h40;
    parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
    parameter [23:0] CLASS_CODE = 24'h000000;
    parameter CMD_INTX_IMPLEMENTED = "TRUE";
    parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
    parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
    parameter [6:0] CRM_MODULE_RSTS = 7'h00;
    parameter [15:0] DEVICE_ID = 16'h0007;
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
    parameter integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
    parameter integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
    parameter integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
    parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
    parameter integer DEV_CAP_RSVD_14_12 = 0;
    parameter integer DEV_CAP_RSVD_17_16 = 0;
    parameter integer DEV_CAP_RSVD_31_29 = 0;
    parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
    parameter DISABLE_ASPM_L1_TIMER = "FALSE";
    parameter DISABLE_BAR_FILTERING = "FALSE";
    parameter DISABLE_ID_CHECK = "FALSE";
    parameter DISABLE_LANE_REVERSAL = "FALSE";
    parameter DISABLE_RX_TC_FILTER = "FALSE";
    parameter DISABLE_SCRAMBLING = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [11:0] DSN_BASE_PTR = 12'h100;
    parameter [15:0] DSN_CAP_ID = 16'h0003;
    parameter [11:0] DSN_CAP_NEXTPTR = 12'h000;
    parameter DSN_CAP_ON = "TRUE";
    parameter [3:0] DSN_CAP_VERSION = 4'h1;
    parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
    parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
    parameter ENTER_RVRY_EI_L0 = "TRUE";
    parameter EXIT_LOOPBACK_ON_EI = "TRUE";
    parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
    parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
    parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
    parameter [7:0] HEADER_TYPE = 8'h00;
    parameter [4:0] INFER_EI = 5'h00;
    parameter [7:0] INTERRUPT_PIN = 8'h01;
    parameter IS_SWITCH = "FALSE";
    parameter [9:0] LAST_CONFIG_DWORD = 10'h042;
    parameter integer LINK_CAP_ASPM_SUPPORT = 1;
    parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
    parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
    parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
    parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
    parameter integer LINK_CAP_RSVD_23_22 = 0;
    parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
    parameter integer LINK_CONTROL_RCB = 0;
    parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
    parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
    parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
    parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
    parameter [7:0] MSIX_BASE_PTR = 8'h9C;
    parameter [7:0] MSIX_CAP_ID = 8'h11;
    parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
    parameter MSIX_CAP_ON = "FALSE";
    parameter integer MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] MSI_BASE_PTR = 8'h48;
    parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
    parameter [7:0] MSI_CAP_ID = 8'h05;
    parameter integer MSI_CAP_MULTIMSGCAP = 0;
    parameter integer MSI_CAP_MULTIMSG_EXTENSION = 0;
    parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
    parameter MSI_CAP_ON = "FALSE";
    parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
    parameter integer N_FTS_COMCLK_GEN1 = 255;
    parameter integer N_FTS_COMCLK_GEN2 = 255;
    parameter integer N_FTS_GEN1 = 255;
    parameter integer N_FTS_GEN2 = 255;
    parameter [7:0] PCIE_BASE_PTR = 8'h60;
    parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
    parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
    parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
    parameter [4:0] PCIE_CAP_INT_MSG_NUM = 5'h00;
    parameter [7:0] PCIE_CAP_NEXTPTR = 8'h00;
    parameter PCIE_CAP_ON = "TRUE";
    parameter integer PCIE_CAP_RSVD_15_14 = 0;
    parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
    parameter integer PCIE_REVISION = 2;
    parameter integer PGL0_LANE = 0;
    parameter integer PGL1_LANE = 1;
    parameter integer PGL2_LANE = 2;
    parameter integer PGL3_LANE = 3;
    parameter integer PGL4_LANE = 4;
    parameter integer PGL5_LANE = 5;
    parameter integer PGL6_LANE = 6;
    parameter integer PGL7_LANE = 7;
    parameter integer PL_AUTO_CONFIG = 0;
    parameter PL_FAST_TRAIN = "FALSE";
    parameter [7:0] PM_BASE_PTR = 8'h40;
    parameter integer PM_CAP_AUXCURRENT = 0;
    parameter PM_CAP_D1SUPPORT = "TRUE";
    parameter PM_CAP_D2SUPPORT = "TRUE";
    parameter PM_CAP_DSI = "FALSE";
    parameter [7:0] PM_CAP_ID = 8'h01;
    parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
    parameter PM_CAP_ON = "TRUE";
    parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
    parameter PM_CAP_PME_CLOCK = "FALSE";
    parameter integer PM_CAP_RSVD_04 = 0;
    parameter integer PM_CAP_VERSION = 3;
    parameter PM_CSR_B2B3 = "FALSE";
    parameter PM_CSR_BPCCEN = "FALSE";
    parameter PM_CSR_NOSOFTRST = "TRUE";
    parameter [7:0] PM_DATA0 = 8'h01;
    parameter [7:0] PM_DATA1 = 8'h01;
    parameter [7:0] PM_DATA2 = 8'h01;
    parameter [7:0] PM_DATA3 = 8'h01;
    parameter [7:0] PM_DATA4 = 8'h01;
    parameter [7:0] PM_DATA5 = 8'h01;
    parameter [7:0] PM_DATA6 = 8'h01;
    parameter [7:0] PM_DATA7 = 8'h01;
    parameter [1:0] PM_DATA_SCALE0 = 2'h1;
    parameter [1:0] PM_DATA_SCALE1 = 2'h1;
    parameter [1:0] PM_DATA_SCALE2 = 2'h1;
    parameter [1:0] PM_DATA_SCALE3 = 2'h1;
    parameter [1:0] PM_DATA_SCALE4 = 2'h1;
    parameter [1:0] PM_DATA_SCALE5 = 2'h1;
    parameter [1:0] PM_DATA_SCALE6 = 2'h1;
    parameter [1:0] PM_DATA_SCALE7 = 2'h1;
    parameter integer RECRC_CHK = 0;
    parameter RECRC_CHK_TRIM = "FALSE";
    parameter [7:0] REVISION_ID = 8'h00;
    parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
    parameter SELECT_DLL_IF = "FALSE";
    parameter SIM_VERSION = "1.0";
    parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
    parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
    parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
    parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
    parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
    parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
    parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
    parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
    parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
    parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
    parameter integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
    parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter [15:0] SUBSYSTEM_ID = 16'h0007;
    parameter [15:0] SUBSYSTEM_VENDOR_ID = 16'h10EE;
    parameter TL_RBYPASS = "FALSE";
    parameter integer TL_RX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_RX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_RX_RAM_WRITE_LATENCY = 0;
    parameter TL_TFC_DISABLE = "FALSE";
    parameter TL_TX_CHECKS_DISABLE = "FALSE";
    parameter integer TL_TX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_TX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_TX_RAM_WRITE_LATENCY = 0;
    parameter UPCONFIG_CAPABLE = "TRUE";
    parameter UPSTREAM_FACING = "TRUE";
    parameter UR_INV_REQ = "TRUE";
    parameter integer USER_CLK_FREQ = 3;
    parameter VC0_CPL_INFINITE = "TRUE";
    parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
    parameter integer VC0_TOTAL_CREDITS_CD = 127;
    parameter integer VC0_TOTAL_CREDITS_CH = 31;
    parameter integer VC0_TOTAL_CREDITS_NPH = 12;
    parameter integer VC0_TOTAL_CREDITS_PD = 288;
    parameter integer VC0_TOTAL_CREDITS_PH = 32;
    parameter integer VC0_TX_LASTPACKET = 31;
    parameter [11:0] VC_BASE_PTR = 12'h10C;
    parameter [15:0] VC_CAP_ID = 16'h0002;
    parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
    parameter VC_CAP_ON = "FALSE";
    parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
    parameter [3:0] VC_CAP_VERSION = 4'h1;
    parameter [15:0] VENDOR_ID = 16'h10EE;
    parameter [11:0] VSEC_BASE_PTR = 12'h160;
    parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
    parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
    parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
    parameter [15:0] VSEC_CAP_ID = 16'h000B;
    parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
    parameter [11:0] VSEC_CAP_NEXTPTR = 12'h000;
    parameter VSEC_CAP_ON = "FALSE";
    parameter [3:0] VSEC_CAP_VERSION = 4'h1;
    output CFGAERECRCCHECKEN;
    output CFGAERECRCGENEN;
    output CFGCOMMANDBUSMASTERENABLE;
    output CFGCOMMANDINTERRUPTDISABLE;
    output CFGCOMMANDIOENABLE;
    output CFGCOMMANDMEMENABLE;
    output CFGCOMMANDSERREN;
    output CFGDEVCONTROL2CPLTIMEOUTDIS;
    output CFGDEVCONTROLAUXPOWEREN;
    output CFGDEVCONTROLCORRERRREPORTINGEN;
    output CFGDEVCONTROLENABLERO;
    output CFGDEVCONTROLEXTTAGEN;
    output CFGDEVCONTROLFATALERRREPORTINGEN;
    output CFGDEVCONTROLNONFATALREPORTINGEN;
    output CFGDEVCONTROLNOSNOOPEN;
    output CFGDEVCONTROLPHANTOMEN;
    output CFGDEVCONTROLURERRREPORTINGEN;
    output CFGDEVSTATUSCORRERRDETECTED;
    output CFGDEVSTATUSFATALERRDETECTED;
    output CFGDEVSTATUSNONFATALERRDETECTED;
    output CFGDEVSTATUSURDETECTED;
    output CFGERRAERHEADERLOGSETN;
    output CFGERRCPLRDYN;
    output CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFM;
    output CFGINTERRUPTRDYN;
    output CFGLINKCONTROLAUTOBANDWIDTHINTEN;
    output CFGLINKCONTROLBANDWIDTHINTEN;
    output CFGLINKCONTROLCLOCKPMEN;
    output CFGLINKCONTROLCOMMONCLOCK;
    output CFGLINKCONTROLEXTENDEDSYNC;
    output CFGLINKCONTROLHWAUTOWIDTHDIS;
    output CFGLINKCONTROLLINKDISABLE;
    output CFGLINKCONTROLRCB;
    output CFGLINKCONTROLRETRAINLINK;
    output CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
    output CFGLINKSTATUSBANDWITHSTATUS;
    output CFGLINKSTATUSDLLACTIVE;
    output CFGLINKSTATUSLINKTRAINING;
    output CFGMSGRECEIVED;
    output CFGMSGRECEIVEDASSERTINTA;
    output CFGMSGRECEIVEDASSERTINTB;
    output CFGMSGRECEIVEDASSERTINTC;
    output CFGMSGRECEIVEDASSERTINTD;
    output CFGMSGRECEIVEDDEASSERTINTA;
    output CFGMSGRECEIVEDDEASSERTINTB;
    output CFGMSGRECEIVEDDEASSERTINTC;
    output CFGMSGRECEIVEDDEASSERTINTD;
    output CFGMSGRECEIVEDERRCOR;
    output CFGMSGRECEIVEDERRFATAL;
    output CFGMSGRECEIVEDERRNONFATAL;
    output CFGMSGRECEIVEDPMASNAK;
    output CFGMSGRECEIVEDPMETO;
    output CFGMSGRECEIVEDPMETOACK;
    output CFGMSGRECEIVEDPMPME;
    output CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
    output CFGMSGRECEIVEDUNLOCK;
    output CFGPMCSRPMEEN;
    output CFGPMCSRPMESTATUS;
    output CFGPMRCVASREQL1N;
    output CFGPMRCVENTERL1N;
    output CFGPMRCVENTERL23N;
    output CFGPMRCVREQACKN;
    output CFGRDWRDONEN;
    output CFGSLOTCONTROLELECTROMECHILCTLPULSE;
    output CFGTRANSACTION;
    output CFGTRANSACTIONTYPE;
    output DBGSCLRA;
    output DBGSCLRB;
    output DBGSCLRC;
    output DBGSCLRD;
    output DBGSCLRE;
    output DBGSCLRF;
    output DBGSCLRG;
    output DBGSCLRH;
    output DBGSCLRI;
    output DBGSCLRJ;
    output DBGSCLRK;
    output DRPDRDY;
    output LL2BADDLLPERRN;
    output LL2BADTLPERRN;
    output LL2PROTOCOLERRN;
    output LL2REPLAYROERRN;
    output LL2REPLAYTOERRN;
    output LL2SUSPENDOKN;
    output LL2TFCINIT1SEQN;
    output LL2TFCINIT2SEQN;
    output LNKCLKEN;
    output MIMRXRCE;
    output MIMRXREN;
    output MIMRXWEN;
    output MIMTXRCE;
    output MIMTXREN;
    output MIMTXWEN;
    output PIPERX0POLARITY;
    output PIPERX1POLARITY;
    output PIPERX2POLARITY;
    output PIPERX3POLARITY;
    output PIPERX4POLARITY;
    output PIPERX5POLARITY;
    output PIPERX6POLARITY;
    output PIPERX7POLARITY;
    output PIPETX0COMPLIANCE;
    output PIPETX0ELECIDLE;
    output PIPETX1COMPLIANCE;
    output PIPETX1ELECIDLE;
    output PIPETX2COMPLIANCE;
    output PIPETX2ELECIDLE;
    output PIPETX3COMPLIANCE;
    output PIPETX3ELECIDLE;
    output PIPETX4COMPLIANCE;
    output PIPETX4ELECIDLE;
    output PIPETX5COMPLIANCE;
    output PIPETX5ELECIDLE;
    output PIPETX6COMPLIANCE;
    output PIPETX6ELECIDLE;
    output PIPETX7COMPLIANCE;
    output PIPETX7ELECIDLE;
    output PIPETXDEEMPH;
    output PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PL2LINKUPN;
    output PL2RECEIVERERRN;
    output PL2RECOVERYN;
    output PL2RXELECIDLE;
    output PL2SUSPENDOK;
    output PLLINKGEN2CAP;
    output PLLINKPARTNERGEN2SUPPORTED;
    output PLLINKUPCFGCAP;
    output PLPHYLNKUPN;
    output PLRECEIVEDHOTRST;
    output PLSELLNKRATE;
    output RECEIVEDFUNCLVLRSTN;
    output TL2ASPMSUSPENDCREDITCHECKOKN;
    output TL2ASPMSUSPENDREQN;
    output TL2PPMSUSPENDOKN;
    output TRNLNKUPN;
    output TRNRDLLPSRCRDYN;
    output TRNRECRCERRN;
    output TRNREOFN;
    output TRNRERRFWDN;
    output TRNRREMN;
    output TRNRSOFN;
    output TRNRSRCDSCN;
    output TRNRSRCRDYN;
    output TRNTCFGREQN;
    output TRNTDLLPDSTRDYN;
    output TRNTDSTRDYN;
    output TRNTERRDROPN;
    output USERRSTN;
    output [11:0] DBGVECC;
    output [11:0] PLDBGVEC;
    output [11:0] TRNFCCPLD;
    output [11:0] TRNFCNPD;
    output [11:0] TRNFCPD;
    output [12:0] MIMRXRADDR;
    output [12:0] MIMRXWADDR;
    output [12:0] MIMTXRADDR;
    output [12:0] MIMTXWADDR;
    output [15:0] CFGMSGDATA;
    output [15:0] DRPDO;
    output [15:0] PIPETX0DATA;
    output [15:0] PIPETX1DATA;
    output [15:0] PIPETX2DATA;
    output [15:0] PIPETX3DATA;
    output [15:0] PIPETX4DATA;
    output [15:0] PIPETX5DATA;
    output [15:0] PIPETX6DATA;
    output [15:0] PIPETX7DATA;
    output [1:0] CFGLINKCONTROLASPMCONTROL;
    output [1:0] CFGLINKSTATUSCURRENTSPEED;
    output [1:0] CFGPMCSRPOWERSTATE;
    output [1:0] PIPETX0CHARISK;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX1CHARISK;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX2CHARISK;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX3CHARISK;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX4CHARISK;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX5CHARISK;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX6CHARISK;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX7CHARISK;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PLLANEREVERSALMODE;
    output [1:0] PLRXPMSTATE;
    output [1:0] PLSELLNKWIDTH;
    output [2:0] CFGDEVCONTROLMAXPAYLOAD;
    output [2:0] CFGDEVCONTROLMAXREADREQ;
    output [2:0] CFGINTERRUPTMMENABLE;
    output [2:0] CFGPCIELINKSTATE;
    output [2:0] PIPETXMARGIN;
    output [2:0] PLINITIALLINKWIDTH;
    output [2:0] PLTXPMSTATE;
    output [31:0] CFGDO;
    output [31:0] TRNRDLLPDATA;
    output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL;
    output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH;
    output [5:0] PLLTSSMSTATE;
    output [5:0] TRNTBUFAV;
    output [63:0] DBGVECA;
    output [63:0] DBGVECB;
    output [63:0] TRNRD;
    output [67:0] MIMRXWDATA;
    output [68:0] MIMTXWDATA;
    output [6:0] CFGTRANSACTIONADDR;
    output [6:0] CFGVCTCVCMAP;
    output [6:0] TRNRBARHITN;
    output [7:0] CFGINTERRUPTDO;
    output [7:0] TRNFCCPLH;
    output [7:0] TRNFCNPH;
    output [7:0] TRNFCPH;
    input CFGERRACSN;
    input CFGERRCORN;
    input CFGERRCPLABORTN;
    input CFGERRCPLTIMEOUTN;
    input CFGERRCPLUNEXPECTN;
    input CFGERRECRCN;
    input CFGERRLOCKEDN;
    input CFGERRPOSTEDN;
    input CFGERRURN;
    input CFGINTERRUPTASSERTN;
    input CFGINTERRUPTN;
    input CFGPMDIRECTASPML1N;
    input CFGPMSENDPMACKN;
    input CFGPMSENDPMETON;
    input CFGPMSENDPMNAKN;
    input CFGPMTURNOFFOKN;
    input CFGPMWAKEN;
    input CFGRDENN;
    input CFGTRNPENDINGN;
    input CFGWRENN;
    input CFGWRREADONLYN;
    input CFGWRRW1CASRWN;
    input CMRSTN;
    input CMSTICKYRSTN;
    input DBGSUBMODE;
    input DLRSTN;
    input DRPCLK;
    input DRPDEN;
    input DRPDWE;
    input FUNCLVLRSTN;
    input LL2SENDASREQL1N;
    input LL2SENDENTERL1N;
    input LL2SENDENTERL23N;
    input LL2SUSPENDNOWN;
    input LL2TLPRCVN;
    input PIPECLK;
    input PIPERX0CHANISALIGNED;
    input PIPERX0ELECIDLE;
    input PIPERX0PHYSTATUS;
    input PIPERX0VALID;
    input PIPERX1CHANISALIGNED;
    input PIPERX1ELECIDLE;
    input PIPERX1PHYSTATUS;
    input PIPERX1VALID;
    input PIPERX2CHANISALIGNED;
    input PIPERX2ELECIDLE;
    input PIPERX2PHYSTATUS;
    input PIPERX2VALID;
    input PIPERX3CHANISALIGNED;
    input PIPERX3ELECIDLE;
    input PIPERX3PHYSTATUS;
    input PIPERX3VALID;
    input PIPERX4CHANISALIGNED;
    input PIPERX4ELECIDLE;
    input PIPERX4PHYSTATUS;
    input PIPERX4VALID;
    input PIPERX5CHANISALIGNED;
    input PIPERX5ELECIDLE;
    input PIPERX5PHYSTATUS;
    input PIPERX5VALID;
    input PIPERX6CHANISALIGNED;
    input PIPERX6ELECIDLE;
    input PIPERX6PHYSTATUS;
    input PIPERX6VALID;
    input PIPERX7CHANISALIGNED;
    input PIPERX7ELECIDLE;
    input PIPERX7PHYSTATUS;
    input PIPERX7VALID;
    input PLDIRECTEDLINKAUTON;
    input PLDIRECTEDLINKSPEED;
    input PLDOWNSTREAMDEEMPHSOURCE;
    input PLRSTN;
    input PLTRANSMITHOTRST;
    input PLUPSTREAMPREFERDEEMPH;
    input SYSRSTN;
    input TL2ASPMSUSPENDCREDITCHECKN;
    input TL2PPMSUSPENDREQN;
    input TLRSTN;
    input TRNRDSTRDYN;
    input TRNRNPOKN;
    input TRNTCFGGNTN;
    input TRNTDLLPSRCRDYN;
    input TRNTECRCGENN;
    input TRNTEOFN;
    input TRNTERRFWDN;
    input TRNTREMN;
    input TRNTSOFN;
    input TRNTSRCDSCN;
    input TRNTSRCRDYN;
    input TRNTSTRN;
    input USERCLK;
    input [127:0] CFGERRAERHEADERLOG;
    input [15:0] DRPDI;
    input [15:0] PIPERX0DATA;
    input [15:0] PIPERX1DATA;
    input [15:0] PIPERX2DATA;
    input [15:0] PIPERX3DATA;
    input [15:0] PIPERX4DATA;
    input [15:0] PIPERX5DATA;
    input [15:0] PIPERX6DATA;
    input [15:0] PIPERX7DATA;
    input [1:0] DBGMODE;
    input [1:0] PIPERX0CHARISK;
    input [1:0] PIPERX1CHARISK;
    input [1:0] PIPERX2CHARISK;
    input [1:0] PIPERX3CHARISK;
    input [1:0] PIPERX4CHARISK;
    input [1:0] PIPERX5CHARISK;
    input [1:0] PIPERX6CHARISK;
    input [1:0] PIPERX7CHARISK;
    input [1:0] PLDIRECTEDLINKCHANGE;
    input [1:0] PLDIRECTEDLINKWIDTH;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [2:0] PIPERX0STATUS;
    input [2:0] PIPERX1STATUS;
    input [2:0] PIPERX2STATUS;
    input [2:0] PIPERX3STATUS;
    input [2:0] PIPERX4STATUS;
    input [2:0] PIPERX5STATUS;
    input [2:0] PIPERX6STATUS;
    input [2:0] PIPERX7STATUS;
    input [2:0] PLDBGMODE;
    input [2:0] TRNFCSEL;
    input [31:0] CFGDI;
    input [31:0] TRNTDLLPDATA;
    input [3:0] CFGBYTEENN;
    input [47:0] CFGERRTLPCPLHEADER;
    input [4:0] CFGDSDEVICENUMBER;
    input [4:0] PL2DIRECTEDLSTATE;
    input [63:0] CFGDSN;
    input [63:0] TRNTD;
    input [67:0] MIMRXRDATA;
    input [68:0] MIMTXRDATA;
    input [7:0] CFGDSBUSNUMBER;
    input [7:0] CFGINTERRUPTDI;
    input [7:0] CFGPORTNUMBER;
    input [8:0] DRPDADDR;
    input [9:0] CFGDWADDR;
endmodule

module PCIE_2_1 (...);
    parameter [11:0] AER_BASE_PTR = 12'h140;
    parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [15:0] AER_CAP_ID = 16'h0001;
    parameter AER_CAP_MULTIHEADER = "FALSE";
    parameter [11:0] AER_CAP_NEXTPTR = 12'h178;
    parameter AER_CAP_ON = "FALSE";
    parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000;
    parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
    parameter [3:0] AER_CAP_VERSION = 4'h2;
    parameter ALLOW_X8_GEN2 = "FALSE";
    parameter [31:0] BAR0 = 32'hFFFFFF00;
    parameter [31:0] BAR1 = 32'hFFFF0000;
    parameter [31:0] BAR2 = 32'hFFFF000C;
    parameter [31:0] BAR3 = 32'hFFFFFFFF;
    parameter [31:0] BAR4 = 32'h00000000;
    parameter [31:0] BAR5 = 32'h00000000;
    parameter [7:0] CAPABILITIES_PTR = 8'h40;
    parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
    parameter integer CFG_ECRC_ERR_CPLSTAT = 0;
    parameter [23:0] CLASS_CODE = 24'h000000;
    parameter CMD_INTX_IMPLEMENTED = "TRUE";
    parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
    parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
    parameter [6:0] CRM_MODULE_RSTS = 7'h00;
    parameter DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE";
    parameter DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE";
    parameter DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE";
    parameter DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE";
    parameter [1:0] DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0;
    parameter DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE";
    parameter [1:0] DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0;
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
    parameter integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
    parameter integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
    parameter integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
    parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
    parameter integer DEV_CAP_RSVD_14_12 = 0;
    parameter integer DEV_CAP_RSVD_17_16 = 0;
    parameter integer DEV_CAP_RSVD_31_29 = 0;
    parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
    parameter DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE";
    parameter DISABLE_ASPM_L1_TIMER = "FALSE";
    parameter DISABLE_BAR_FILTERING = "FALSE";
    parameter DISABLE_ERR_MSG = "FALSE";
    parameter DISABLE_ID_CHECK = "FALSE";
    parameter DISABLE_LANE_REVERSAL = "FALSE";
    parameter DISABLE_LOCKED_FILTER = "FALSE";
    parameter DISABLE_PPM_FILTER = "FALSE";
    parameter DISABLE_RX_POISONED_RESP = "FALSE";
    parameter DISABLE_RX_TC_FILTER = "FALSE";
    parameter DISABLE_SCRAMBLING = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [11:0] DSN_BASE_PTR = 12'h100;
    parameter [15:0] DSN_CAP_ID = 16'h0003;
    parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C;
    parameter DSN_CAP_ON = "TRUE";
    parameter [3:0] DSN_CAP_VERSION = 4'h1;
    parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
    parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
    parameter ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE";
    parameter ENTER_RVRY_EI_L0 = "TRUE";
    parameter EXIT_LOOPBACK_ON_EI = "TRUE";
    parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
    parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
    parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
    parameter [7:0] HEADER_TYPE = 8'h00;
    parameter [4:0] INFER_EI = 5'h00;
    parameter [7:0] INTERRUPT_PIN = 8'h01;
    parameter INTERRUPT_STAT_AUTO = "TRUE";
    parameter IS_SWITCH = "FALSE";
    parameter [9:0] LAST_CONFIG_DWORD = 10'h3FF;
    parameter LINK_CAP_ASPM_OPTIONALITY = "TRUE";
    parameter integer LINK_CAP_ASPM_SUPPORT = 1;
    parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
    parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
    parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
    parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
    parameter integer LINK_CAP_RSVD_23 = 0;
    parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
    parameter integer LINK_CONTROL_RCB = 0;
    parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
    parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
    parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
    parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
    parameter MPS_FORCE = "FALSE";
    parameter [7:0] MSIX_BASE_PTR = 8'h9C;
    parameter [7:0] MSIX_CAP_ID = 8'h11;
    parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
    parameter MSIX_CAP_ON = "FALSE";
    parameter integer MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] MSI_BASE_PTR = 8'h48;
    parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
    parameter [7:0] MSI_CAP_ID = 8'h05;
    parameter integer MSI_CAP_MULTIMSGCAP = 0;
    parameter integer MSI_CAP_MULTIMSG_EXTENSION = 0;
    parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
    parameter MSI_CAP_ON = "FALSE";
    parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
    parameter integer N_FTS_COMCLK_GEN1 = 255;
    parameter integer N_FTS_COMCLK_GEN2 = 255;
    parameter integer N_FTS_GEN1 = 255;
    parameter integer N_FTS_GEN2 = 255;
    parameter [7:0] PCIE_BASE_PTR = 8'h60;
    parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
    parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
    parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
    parameter [7:0] PCIE_CAP_NEXTPTR = 8'h9C;
    parameter PCIE_CAP_ON = "TRUE";
    parameter integer PCIE_CAP_RSVD_15_14 = 0;
    parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
    parameter integer PCIE_REVISION = 2;
    parameter integer PL_AUTO_CONFIG = 0;
    parameter PL_FAST_TRAIN = "FALSE";
    parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000;
    parameter PM_ASPML0S_TIMEOUT_EN = "FALSE";
    parameter integer PM_ASPML0S_TIMEOUT_FUNC = 0;
    parameter PM_ASPM_FASTEXIT = "FALSE";
    parameter [7:0] PM_BASE_PTR = 8'h40;
    parameter integer PM_CAP_AUXCURRENT = 0;
    parameter PM_CAP_D1SUPPORT = "TRUE";
    parameter PM_CAP_D2SUPPORT = "TRUE";
    parameter PM_CAP_DSI = "FALSE";
    parameter [7:0] PM_CAP_ID = 8'h01;
    parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
    parameter PM_CAP_ON = "TRUE";
    parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
    parameter PM_CAP_PME_CLOCK = "FALSE";
    parameter integer PM_CAP_RSVD_04 = 0;
    parameter integer PM_CAP_VERSION = 3;
    parameter PM_CSR_B2B3 = "FALSE";
    parameter PM_CSR_BPCCEN = "FALSE";
    parameter PM_CSR_NOSOFTRST = "TRUE";
    parameter [7:0] PM_DATA0 = 8'h01;
    parameter [7:0] PM_DATA1 = 8'h01;
    parameter [7:0] PM_DATA2 = 8'h01;
    parameter [7:0] PM_DATA3 = 8'h01;
    parameter [7:0] PM_DATA4 = 8'h01;
    parameter [7:0] PM_DATA5 = 8'h01;
    parameter [7:0] PM_DATA6 = 8'h01;
    parameter [7:0] PM_DATA7 = 8'h01;
    parameter [1:0] PM_DATA_SCALE0 = 2'h1;
    parameter [1:0] PM_DATA_SCALE1 = 2'h1;
    parameter [1:0] PM_DATA_SCALE2 = 2'h1;
    parameter [1:0] PM_DATA_SCALE3 = 2'h1;
    parameter [1:0] PM_DATA_SCALE4 = 2'h1;
    parameter [1:0] PM_DATA_SCALE5 = 2'h1;
    parameter [1:0] PM_DATA_SCALE6 = 2'h1;
    parameter [1:0] PM_DATA_SCALE7 = 2'h1;
    parameter PM_MF = "FALSE";
    parameter [11:0] RBAR_BASE_PTR = 12'h178;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00;
    parameter [15:0] RBAR_CAP_ID = 16'h0015;
    parameter [2:0] RBAR_CAP_INDEX0 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX1 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX2 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX3 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX4 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX5 = 3'h0;
    parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000;
    parameter RBAR_CAP_ON = "FALSE";
    parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000;
    parameter [3:0] RBAR_CAP_VERSION = 4'h1;
    parameter [2:0] RBAR_NUM = 3'h1;
    parameter integer RECRC_CHK = 0;
    parameter RECRC_CHK_TRIM = "FALSE";
    parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
    parameter [1:0] RP_AUTO_SPD = 2'h1;
    parameter [4:0] RP_AUTO_SPD_LOOPCNT = 5'h1F;
    parameter SELECT_DLL_IF = "FALSE";
    parameter SIM_VERSION = "1.0";
    parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
    parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
    parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
    parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
    parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
    parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
    parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
    parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
    parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
    parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
    parameter integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
    parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SSL_MESSAGE_AUTO = "FALSE";
    parameter TECRC_EP_INV = "FALSE";
    parameter TL_RBYPASS = "FALSE";
    parameter integer TL_RX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_RX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_RX_RAM_WRITE_LATENCY = 0;
    parameter TL_TFC_DISABLE = "FALSE";
    parameter TL_TX_CHECKS_DISABLE = "FALSE";
    parameter integer TL_TX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_TX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_TX_RAM_WRITE_LATENCY = 0;
    parameter TRN_DW = "FALSE";
    parameter TRN_NP_FC = "FALSE";
    parameter UPCONFIG_CAPABLE = "TRUE";
    parameter UPSTREAM_FACING = "TRUE";
    parameter UR_ATOMIC = "TRUE";
    parameter UR_CFG1 = "TRUE";
    parameter UR_INV_REQ = "TRUE";
    parameter UR_PRS_RESPONSE = "TRUE";
    parameter USER_CLK2_DIV2 = "FALSE";
    parameter integer USER_CLK_FREQ = 3;
    parameter USE_RID_PINS = "FALSE";
    parameter VC0_CPL_INFINITE = "TRUE";
    parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
    parameter integer VC0_TOTAL_CREDITS_CD = 127;
    parameter integer VC0_TOTAL_CREDITS_CH = 31;
    parameter integer VC0_TOTAL_CREDITS_NPD = 24;
    parameter integer VC0_TOTAL_CREDITS_NPH = 12;
    parameter integer VC0_TOTAL_CREDITS_PD = 288;
    parameter integer VC0_TOTAL_CREDITS_PH = 32;
    parameter integer VC0_TX_LASTPACKET = 31;
    parameter [11:0] VC_BASE_PTR = 12'h10C;
    parameter [15:0] VC_CAP_ID = 16'h0002;
    parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
    parameter VC_CAP_ON = "FALSE";
    parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
    parameter [3:0] VC_CAP_VERSION = 4'h1;
    parameter [11:0] VSEC_BASE_PTR = 12'h128;
    parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
    parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
    parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
    parameter [15:0] VSEC_CAP_ID = 16'h000B;
    parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
    parameter [11:0] VSEC_CAP_NEXTPTR = 12'h140;
    parameter VSEC_CAP_ON = "FALSE";
    parameter [3:0] VSEC_CAP_VERSION = 4'h1;
    output CFGAERECRCCHECKEN;
    output CFGAERECRCGENEN;
    output CFGAERROOTERRCORRERRRECEIVED;
    output CFGAERROOTERRCORRERRREPORTINGEN;
    output CFGAERROOTERRFATALERRRECEIVED;
    output CFGAERROOTERRFATALERRREPORTINGEN;
    output CFGAERROOTERRNONFATALERRRECEIVED;
    output CFGAERROOTERRNONFATALERRREPORTINGEN;
    output CFGBRIDGESERREN;
    output CFGCOMMANDBUSMASTERENABLE;
    output CFGCOMMANDINTERRUPTDISABLE;
    output CFGCOMMANDIOENABLE;
    output CFGCOMMANDMEMENABLE;
    output CFGCOMMANDSERREN;
    output CFGDEVCONTROL2ARIFORWARDEN;
    output CFGDEVCONTROL2ATOMICEGRESSBLOCK;
    output CFGDEVCONTROL2ATOMICREQUESTEREN;
    output CFGDEVCONTROL2CPLTIMEOUTDIS;
    output CFGDEVCONTROL2IDOCPLEN;
    output CFGDEVCONTROL2IDOREQEN;
    output CFGDEVCONTROL2LTREN;
    output CFGDEVCONTROL2TLPPREFIXBLOCK;
    output CFGDEVCONTROLAUXPOWEREN;
    output CFGDEVCONTROLCORRERRREPORTINGEN;
    output CFGDEVCONTROLENABLERO;
    output CFGDEVCONTROLEXTTAGEN;
    output CFGDEVCONTROLFATALERRREPORTINGEN;
    output CFGDEVCONTROLNONFATALREPORTINGEN;
    output CFGDEVCONTROLNOSNOOPEN;
    output CFGDEVCONTROLPHANTOMEN;
    output CFGDEVCONTROLURERRREPORTINGEN;
    output CFGDEVSTATUSCORRERRDETECTED;
    output CFGDEVSTATUSFATALERRDETECTED;
    output CFGDEVSTATUSNONFATALERRDETECTED;
    output CFGDEVSTATUSURDETECTED;
    output CFGERRAERHEADERLOGSETN;
    output CFGERRCPLRDYN;
    output CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFM;
    output CFGINTERRUPTRDYN;
    output CFGLINKCONTROLAUTOBANDWIDTHINTEN;
    output CFGLINKCONTROLBANDWIDTHINTEN;
    output CFGLINKCONTROLCLOCKPMEN;
    output CFGLINKCONTROLCOMMONCLOCK;
    output CFGLINKCONTROLEXTENDEDSYNC;
    output CFGLINKCONTROLHWAUTOWIDTHDIS;
    output CFGLINKCONTROLLINKDISABLE;
    output CFGLINKCONTROLRCB;
    output CFGLINKCONTROLRETRAINLINK;
    output CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
    output CFGLINKSTATUSBANDWIDTHSTATUS;
    output CFGLINKSTATUSDLLACTIVE;
    output CFGLINKSTATUSLINKTRAINING;
    output CFGMGMTRDWRDONEN;
    output CFGMSGRECEIVED;
    output CFGMSGRECEIVEDASSERTINTA;
    output CFGMSGRECEIVEDASSERTINTB;
    output CFGMSGRECEIVEDASSERTINTC;
    output CFGMSGRECEIVEDASSERTINTD;
    output CFGMSGRECEIVEDDEASSERTINTA;
    output CFGMSGRECEIVEDDEASSERTINTB;
    output CFGMSGRECEIVEDDEASSERTINTC;
    output CFGMSGRECEIVEDDEASSERTINTD;
    output CFGMSGRECEIVEDERRCOR;
    output CFGMSGRECEIVEDERRFATAL;
    output CFGMSGRECEIVEDERRNONFATAL;
    output CFGMSGRECEIVEDPMASNAK;
    output CFGMSGRECEIVEDPMETO;
    output CFGMSGRECEIVEDPMETOACK;
    output CFGMSGRECEIVEDPMPME;
    output CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
    output CFGMSGRECEIVEDUNLOCK;
    output CFGPMCSRPMEEN;
    output CFGPMCSRPMESTATUS;
    output CFGPMRCVASREQL1N;
    output CFGPMRCVENTERL1N;
    output CFGPMRCVENTERL23N;
    output CFGPMRCVREQACKN;
    output CFGROOTCONTROLPMEINTEN;
    output CFGROOTCONTROLSYSERRCORRERREN;
    output CFGROOTCONTROLSYSERRFATALERREN;
    output CFGROOTCONTROLSYSERRNONFATALERREN;
    output CFGSLOTCONTROLELECTROMECHILCTLPULSE;
    output CFGTRANSACTION;
    output CFGTRANSACTIONTYPE;
    output DBGSCLRA;
    output DBGSCLRB;
    output DBGSCLRC;
    output DBGSCLRD;
    output DBGSCLRE;
    output DBGSCLRF;
    output DBGSCLRG;
    output DBGSCLRH;
    output DBGSCLRI;
    output DBGSCLRJ;
    output DBGSCLRK;
    output DRPRDY;
    output LL2BADDLLPERR;
    output LL2BADTLPERR;
    output LL2PROTOCOLERR;
    output LL2RECEIVERERR;
    output LL2REPLAYROERR;
    output LL2REPLAYTOERR;
    output LL2SUSPENDOK;
    output LL2TFCINIT1SEQ;
    output LL2TFCINIT2SEQ;
    output LL2TXIDLE;
    output LNKCLKEN;
    output MIMRXREN;
    output MIMRXWEN;
    output MIMTXREN;
    output MIMTXWEN;
    output PIPERX0POLARITY;
    output PIPERX1POLARITY;
    output PIPERX2POLARITY;
    output PIPERX3POLARITY;
    output PIPERX4POLARITY;
    output PIPERX5POLARITY;
    output PIPERX6POLARITY;
    output PIPERX7POLARITY;
    output PIPETX0COMPLIANCE;
    output PIPETX0ELECIDLE;
    output PIPETX1COMPLIANCE;
    output PIPETX1ELECIDLE;
    output PIPETX2COMPLIANCE;
    output PIPETX2ELECIDLE;
    output PIPETX3COMPLIANCE;
    output PIPETX3ELECIDLE;
    output PIPETX4COMPLIANCE;
    output PIPETX4ELECIDLE;
    output PIPETX5COMPLIANCE;
    output PIPETX5ELECIDLE;
    output PIPETX6COMPLIANCE;
    output PIPETX6ELECIDLE;
    output PIPETX7COMPLIANCE;
    output PIPETX7ELECIDLE;
    output PIPETXDEEMPH;
    output PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PL2L0REQ;
    output PL2LINKUP;
    output PL2RECEIVERERR;
    output PL2RECOVERY;
    output PL2RXELECIDLE;
    output PL2SUSPENDOK;
    output PLDIRECTEDCHANGEDONE;
    output PLLINKGEN2CAP;
    output PLLINKPARTNERGEN2SUPPORTED;
    output PLLINKUPCFGCAP;
    output PLPHYLNKUPN;
    output PLRECEIVEDHOTRST;
    output PLSELLNKRATE;
    output RECEIVEDFUNCLVLRSTN;
    output TL2ASPMSUSPENDCREDITCHECKOK;
    output TL2ASPMSUSPENDREQ;
    output TL2ERRFCPE;
    output TL2ERRMALFORMED;
    output TL2ERRRXOVERFLOW;
    output TL2PPMSUSPENDOK;
    output TRNLNKUP;
    output TRNRECRCERR;
    output TRNREOF;
    output TRNRERRFWD;
    output TRNRSOF;
    output TRNRSRCDSC;
    output TRNRSRCRDY;
    output TRNTCFGREQ;
    output TRNTDLLPDSTRDY;
    output TRNTERRDROP;
    output USERRSTN;
    output [11:0] DBGVECC;
    output [11:0] PLDBGVEC;
    output [11:0] TRNFCCPLD;
    output [11:0] TRNFCNPD;
    output [11:0] TRNFCPD;
    output [127:0] TRNRD;
    output [12:0] MIMRXRADDR;
    output [12:0] MIMRXWADDR;
    output [12:0] MIMTXRADDR;
    output [12:0] MIMTXWADDR;
    output [15:0] CFGMSGDATA;
    output [15:0] DRPDO;
    output [15:0] PIPETX0DATA;
    output [15:0] PIPETX1DATA;
    output [15:0] PIPETX2DATA;
    output [15:0] PIPETX3DATA;
    output [15:0] PIPETX4DATA;
    output [15:0] PIPETX5DATA;
    output [15:0] PIPETX6DATA;
    output [15:0] PIPETX7DATA;
    output [1:0] CFGLINKCONTROLASPMCONTROL;
    output [1:0] CFGLINKSTATUSCURRENTSPEED;
    output [1:0] CFGPMCSRPOWERSTATE;
    output [1:0] PIPETX0CHARISK;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX1CHARISK;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX2CHARISK;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX3CHARISK;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX4CHARISK;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX5CHARISK;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX6CHARISK;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX7CHARISK;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PL2RXPMSTATE;
    output [1:0] PLLANEREVERSALMODE;
    output [1:0] PLRXPMSTATE;
    output [1:0] PLSELLNKWIDTH;
    output [1:0] TRNRDLLPSRCRDY;
    output [1:0] TRNRREM;
    output [2:0] CFGDEVCONTROLMAXPAYLOAD;
    output [2:0] CFGDEVCONTROLMAXREADREQ;
    output [2:0] CFGINTERRUPTMMENABLE;
    output [2:0] CFGPCIELINKSTATE;
    output [2:0] PIPETXMARGIN;
    output [2:0] PLINITIALLINKWIDTH;
    output [2:0] PLTXPMSTATE;
    output [31:0] CFGMGMTDO;
    output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL;
    output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH;
    output [3:0] TRNTDSTRDY;
    output [4:0] LL2LINKSTATUS;
    output [5:0] PLLTSSMSTATE;
    output [5:0] TRNTBUFAV;
    output [63:0] DBGVECA;
    output [63:0] DBGVECB;
    output [63:0] TL2ERRHDR;
    output [63:0] TRNRDLLPDATA;
    output [67:0] MIMRXWDATA;
    output [68:0] MIMTXWDATA;
    output [6:0] CFGTRANSACTIONADDR;
    output [6:0] CFGVCTCVCMAP;
    output [7:0] CFGINTERRUPTDO;
    output [7:0] TRNFCCPLH;
    output [7:0] TRNFCNPH;
    output [7:0] TRNFCPH;
    output [7:0] TRNRBARHIT;
    input CFGERRACSN;
    input CFGERRATOMICEGRESSBLOCKEDN;
    input CFGERRCORN;
    input CFGERRCPLABORTN;
    input CFGERRCPLTIMEOUTN;
    input CFGERRCPLUNEXPECTN;
    input CFGERRECRCN;
    input CFGERRINTERNALCORN;
    input CFGERRINTERNALUNCORN;
    input CFGERRLOCKEDN;
    input CFGERRMALFORMEDN;
    input CFGERRMCBLOCKEDN;
    input CFGERRNORECOVERYN;
    input CFGERRPOISONEDN;
    input CFGERRPOSTEDN;
    input CFGERRURN;
    input CFGFORCECOMMONCLOCKOFF;
    input CFGFORCEEXTENDEDSYNCON;
    input CFGINTERRUPTASSERTN;
    input CFGINTERRUPTN;
    input CFGINTERRUPTSTATN;
    input CFGMGMTRDENN;
    input CFGMGMTWRENN;
    input CFGMGMTWRREADONLYN;
    input CFGMGMTWRRW1CASRWN;
    input CFGPMFORCESTATEENN;
    input CFGPMHALTASPML0SN;
    input CFGPMHALTASPML1N;
    input CFGPMSENDPMETON;
    input CFGPMTURNOFFOKN;
    input CFGPMWAKEN;
    input CFGTRNPENDINGN;
    input CMRSTN;
    input CMSTICKYRSTN;
    input DBGSUBMODE;
    input DLRSTN;
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input FUNCLVLRSTN;
    input LL2SENDASREQL1;
    input LL2SENDENTERL1;
    input LL2SENDENTERL23;
    input LL2SENDPMACK;
    input LL2SUSPENDNOW;
    input LL2TLPRCV;
    input PIPECLK;
    input PIPERX0CHANISALIGNED;
    input PIPERX0ELECIDLE;
    input PIPERX0PHYSTATUS;
    input PIPERX0VALID;
    input PIPERX1CHANISALIGNED;
    input PIPERX1ELECIDLE;
    input PIPERX1PHYSTATUS;
    input PIPERX1VALID;
    input PIPERX2CHANISALIGNED;
    input PIPERX2ELECIDLE;
    input PIPERX2PHYSTATUS;
    input PIPERX2VALID;
    input PIPERX3CHANISALIGNED;
    input PIPERX3ELECIDLE;
    input PIPERX3PHYSTATUS;
    input PIPERX3VALID;
    input PIPERX4CHANISALIGNED;
    input PIPERX4ELECIDLE;
    input PIPERX4PHYSTATUS;
    input PIPERX4VALID;
    input PIPERX5CHANISALIGNED;
    input PIPERX5ELECIDLE;
    input PIPERX5PHYSTATUS;
    input PIPERX5VALID;
    input PIPERX6CHANISALIGNED;
    input PIPERX6ELECIDLE;
    input PIPERX6PHYSTATUS;
    input PIPERX6VALID;
    input PIPERX7CHANISALIGNED;
    input PIPERX7ELECIDLE;
    input PIPERX7PHYSTATUS;
    input PIPERX7VALID;
    input PLDIRECTEDLINKAUTON;
    input PLDIRECTEDLINKSPEED;
    input PLDIRECTEDLTSSMNEWVLD;
    input PLDIRECTEDLTSSMSTALL;
    input PLDOWNSTREAMDEEMPHSOURCE;
    input PLRSTN;
    input PLTRANSMITHOTRST;
    input PLUPSTREAMPREFERDEEMPH;
    input SYSRSTN;
    input TL2ASPMSUSPENDCREDITCHECK;
    input TL2PPMSUSPENDREQ;
    input TLRSTN;
    input TRNRDSTRDY;
    input TRNRFCPRET;
    input TRNRNPOK;
    input TRNRNPREQ;
    input TRNTCFGGNT;
    input TRNTDLLPSRCRDY;
    input TRNTECRCGEN;
    input TRNTEOF;
    input TRNTERRFWD;
    input TRNTSOF;
    input TRNTSRCDSC;
    input TRNTSRCRDY;
    input TRNTSTR;
    input USERCLK2;
    input USERCLK;
    input [127:0] CFGERRAERHEADERLOG;
    input [127:0] TRNTD;
    input [15:0] CFGDEVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [15:0] CFGVENDID;
    input [15:0] DRPDI;
    input [15:0] PIPERX0DATA;
    input [15:0] PIPERX1DATA;
    input [15:0] PIPERX2DATA;
    input [15:0] PIPERX3DATA;
    input [15:0] PIPERX4DATA;
    input [15:0] PIPERX5DATA;
    input [15:0] PIPERX6DATA;
    input [15:0] PIPERX7DATA;
    input [1:0] CFGPMFORCESTATE;
    input [1:0] DBGMODE;
    input [1:0] PIPERX0CHARISK;
    input [1:0] PIPERX1CHARISK;
    input [1:0] PIPERX2CHARISK;
    input [1:0] PIPERX3CHARISK;
    input [1:0] PIPERX4CHARISK;
    input [1:0] PIPERX5CHARISK;
    input [1:0] PIPERX6CHARISK;
    input [1:0] PIPERX7CHARISK;
    input [1:0] PLDIRECTEDLINKCHANGE;
    input [1:0] PLDIRECTEDLINKWIDTH;
    input [1:0] TRNTREM;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [2:0] CFGFORCEMPS;
    input [2:0] PIPERX0STATUS;
    input [2:0] PIPERX1STATUS;
    input [2:0] PIPERX2STATUS;
    input [2:0] PIPERX3STATUS;
    input [2:0] PIPERX4STATUS;
    input [2:0] PIPERX5STATUS;
    input [2:0] PIPERX6STATUS;
    input [2:0] PIPERX7STATUS;
    input [2:0] PLDBGMODE;
    input [2:0] TRNFCSEL;
    input [31:0] CFGMGMTDI;
    input [31:0] TRNTDLLPDATA;
    input [3:0] CFGMGMTBYTEENN;
    input [47:0] CFGERRTLPCPLHEADER;
    input [4:0] CFGAERINTERRUPTMSGNUM;
    input [4:0] CFGDSDEVICENUMBER;
    input [4:0] CFGPCIECAPINTERRUPTMSGNUM;
    input [4:0] PL2DIRECTEDLSTATE;
    input [5:0] PLDIRECTEDLTSSMNEW;
    input [63:0] CFGDSN;
    input [67:0] MIMRXRDATA;
    input [68:0] MIMTXRDATA;
    input [7:0] CFGDSBUSNUMBER;
    input [7:0] CFGINTERRUPTDI;
    input [7:0] CFGPORTNUMBER;
    input [7:0] CFGREVID;
    input [8:0] DRPADDR;
    input [9:0] CFGMGMTDWADDR;
endmodule

module PCIE_3_0 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
    parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [1:0] GEN3_PCS_AUTO_REALIGN = 2'h1;
    parameter GEN3_PCS_RX_ELECIDLE_INTERNAL = "TRUE";
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [4:0] PF0_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_BIST_REGISTER = 8'h00;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter [15:0] PF0_DEVICE_ID = 16'h0000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
    parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF0_PB_CAP_VER = 4'h1;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter PF0_RBAR_CAP_ENABLE = "FALSE";
    parameter [2:0] PF0_RBAR_CAP_INDEX0 = 3'h0;
    parameter [2:0] PF0_RBAR_CAP_INDEX1 = 3'h0;
    parameter [2:0] PF0_RBAR_CAP_INDEX2 = 3'h0;
    parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF0_RBAR_NUM = 3'h1;
    parameter [7:0] PF0_REVISION_ID = 8'h00;
    parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [4:0] PF1_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_BIST_REGISTER = 8'h00;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [15:0] PF1_DEVICE_ID = 16'h0000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
    parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF1_PB_CAP_VER = 4'h1;
    parameter [7:0] PF1_PM_CAP_ID = 8'h01;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
    parameter PF1_RBAR_CAP_ENABLE = "FALSE";
    parameter [2:0] PF1_RBAR_CAP_INDEX0 = 3'h0;
    parameter [2:0] PF1_RBAR_CAP_INDEX1 = 3'h0;
    parameter [2:0] PF1_RBAR_CAP_INDEX2 = 3'h0;
    parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF1_RBAR_NUM = 3'h1;
    parameter [7:0] PF1_REVISION_ID = 8'h00;
    parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
    parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF1_TPHR_CAP_ENABLE = "FALSE";
    parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_SCRAMBLING = "FALSE";
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
    parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
    parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
    parameter integer PL_N_FTS_GEN1 = 255;
    parameter integer PL_N_FTS_GEN2 = 255;
    parameter integer PL_N_FTS_GEN3 = 255;
    parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
    parameter SIM_VERSION = "1.0";
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SRIOV_CAP_ENABLE = "FALSE";
    parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h0000000;
    parameter [11:0] TL_CREDITS_CD = 12'h3E0;
    parameter [7:0] TL_CREDITS_CH = 8'h20;
    parameter [11:0] TL_CREDITS_NPD = 12'h028;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h198;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
    parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_MODE_ENABLE = "FALSE";
    parameter TL_PF_ENABLE_REG = "FALSE";
    parameter TL_TAG_MGMT_ENABLE = "TRUE";
    parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
    parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF0_PM_CAP_ID = 8'h01;
    parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
    parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF0_TPHR_CAP_ENABLE = "FALSE";
    parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF1_PM_CAP_ID = 8'h01;
    parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
    parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF1_TPHR_CAP_ENABLE = "FALSE";
    parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF2_PM_CAP_ID = 8'h01;
    parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
    parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF2_TPHR_CAP_ENABLE = "FALSE";
    parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF3_PM_CAP_ID = 8'h01;
    parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
    parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF3_TPHR_CAP_ENABLE = "FALSE";
    parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF4_PM_CAP_ID = 8'h01;
    parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
    parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF4_TPHR_CAP_ENABLE = "FALSE";
    parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF5_PM_CAP_ID = 8'h01;
    parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
    parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF5_TPHR_CAP_ENABLE = "FALSE";
    parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output CFGEXTREADRECEIVED;
    output CFGEXTWRITERECEIVED;
    output CFGHOTRESETOUT;
    output CFGINPUTUPDATEDONE;
    output CFGINTERRUPTAOUTPUT;
    output CFGINTERRUPTBOUTPUT;
    output CFGINTERRUPTCOUTPUT;
    output CFGINTERRUPTDOUTPUT;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output CFGINTERRUPTMSISENT;
    output CFGINTERRUPTMSIXFAIL;
    output CFGINTERRUPTMSIXSENT;
    output CFGINTERRUPTSENT;
    output CFGLOCALERROR;
    output CFGLTRENABLE;
    output CFGMCUPDATEDONE;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output CFGMSGTRANSMITDONE;
    output CFGPERFUNCTIONUPDATEDONE;
    output CFGPHYLINKDOWN;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output CFGTPHSTTREADENABLE;
    output CFGTPHSTTWRITEENABLE;
    output DRPRDY;
    output MAXISCQTLAST;
    output MAXISCQTVALID;
    output MAXISRCTLAST;
    output MAXISRCTVALID;
    output PCIERQSEQNUMVLD;
    output PCIERQTAGVLD;
    output PIPERX0POLARITY;
    output PIPERX1POLARITY;
    output PIPERX2POLARITY;
    output PIPERX3POLARITY;
    output PIPERX4POLARITY;
    output PIPERX5POLARITY;
    output PIPERX6POLARITY;
    output PIPERX7POLARITY;
    output PIPETX0COMPLIANCE;
    output PIPETX0DATAVALID;
    output PIPETX0ELECIDLE;
    output PIPETX0STARTBLOCK;
    output PIPETX1COMPLIANCE;
    output PIPETX1DATAVALID;
    output PIPETX1ELECIDLE;
    output PIPETX1STARTBLOCK;
    output PIPETX2COMPLIANCE;
    output PIPETX2DATAVALID;
    output PIPETX2ELECIDLE;
    output PIPETX2STARTBLOCK;
    output PIPETX3COMPLIANCE;
    output PIPETX3DATAVALID;
    output PIPETX3ELECIDLE;
    output PIPETX3STARTBLOCK;
    output PIPETX4COMPLIANCE;
    output PIPETX4DATAVALID;
    output PIPETX4ELECIDLE;
    output PIPETX4STARTBLOCK;
    output PIPETX5COMPLIANCE;
    output PIPETX5DATAVALID;
    output PIPETX5ELECIDLE;
    output PIPETX5STARTBLOCK;
    output PIPETX6COMPLIANCE;
    output PIPETX6DATAVALID;
    output PIPETX6ELECIDLE;
    output PIPETX6STARTBLOCK;
    output PIPETX7COMPLIANCE;
    output PIPETX7DATAVALID;
    output PIPETX7ELECIDLE;
    output PIPETX7STARTBLOCK;
    output PIPETXDEEMPH;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PIPETXSWING;
    output PLEQINPROGRESS;
    output [11:0] CFGFCCPLD;
    output [11:0] CFGFCNPD;
    output [11:0] CFGFCPD;
    output [11:0] CFGVFSTATUS;
    output [143:0] MIREPLAYRAMWRITEDATA;
    output [143:0] MIREQUESTRAMWRITEDATA;
    output [15:0] CFGPERFUNCSTATUSDATA;
    output [15:0] DBGDATAOUT;
    output [15:0] DRPDO;
    output [17:0] CFGVFPOWERSTATE;
    output [17:0] CFGVFTPHSTMODE;
    output [1:0] CFGDPASUBSTATECHANGE;
    output [1:0] CFGFLRINPROCESS;
    output [1:0] CFGINTERRUPTMSIENABLE;
    output [1:0] CFGINTERRUPTMSIXENABLE;
    output [1:0] CFGINTERRUPTMSIXMASK;
    output [1:0] CFGLINKPOWERSTATE;
    output [1:0] CFGOBFFENABLE;
    output [1:0] CFGPHYLINKSTATUS;
    output [1:0] CFGRCBSTATUS;
    output [1:0] CFGTPHREQUESTERENABLE;
    output [1:0] MIREPLAYRAMREADENABLE;
    output [1:0] MIREPLAYRAMWRITEENABLE;
    output [1:0] PCIERQTAGAV;
    output [1:0] PCIETFCNPDAV;
    output [1:0] PCIETFCNPHAV;
    output [1:0] PIPERX0EQCONTROL;
    output [1:0] PIPERX1EQCONTROL;
    output [1:0] PIPERX2EQCONTROL;
    output [1:0] PIPERX3EQCONTROL;
    output [1:0] PIPERX4EQCONTROL;
    output [1:0] PIPERX5EQCONTROL;
    output [1:0] PIPERX6EQCONTROL;
    output [1:0] PIPERX7EQCONTROL;
    output [1:0] PIPETX0CHARISK;
    output [1:0] PIPETX0EQCONTROL;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX0SYNCHEADER;
    output [1:0] PIPETX1CHARISK;
    output [1:0] PIPETX1EQCONTROL;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX1SYNCHEADER;
    output [1:0] PIPETX2CHARISK;
    output [1:0] PIPETX2EQCONTROL;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX2SYNCHEADER;
    output [1:0] PIPETX3CHARISK;
    output [1:0] PIPETX3EQCONTROL;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX3SYNCHEADER;
    output [1:0] PIPETX4CHARISK;
    output [1:0] PIPETX4EQCONTROL;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX4SYNCHEADER;
    output [1:0] PIPETX5CHARISK;
    output [1:0] PIPETX5EQCONTROL;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX5SYNCHEADER;
    output [1:0] PIPETX6CHARISK;
    output [1:0] PIPETX6EQCONTROL;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX6SYNCHEADER;
    output [1:0] PIPETX7CHARISK;
    output [1:0] PIPETX7EQCONTROL;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PIPETX7SYNCHEADER;
    output [1:0] PIPETXRATE;
    output [1:0] PLEQPHASE;
    output [255:0] MAXISCQTDATA;
    output [255:0] MAXISRCTDATA;
    output [2:0] CFGCURRENTSPEED;
    output [2:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [2:0] CFGTPHFUNCTIONNUM;
    output [2:0] PIPERX0EQPRESET;
    output [2:0] PIPERX1EQPRESET;
    output [2:0] PIPERX2EQPRESET;
    output [2:0] PIPERX3EQPRESET;
    output [2:0] PIPERX4EQPRESET;
    output [2:0] PIPERX5EQPRESET;
    output [2:0] PIPERX6EQPRESET;
    output [2:0] PIPERX7EQPRESET;
    output [2:0] PIPETXMARGIN;
    output [31:0] CFGEXTWRITEDATA;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [31:0] CFGMGMTREADDATA;
    output [31:0] CFGTPHSTTWRITEDATA;
    output [31:0] PIPETX0DATA;
    output [31:0] PIPETX1DATA;
    output [31:0] PIPETX2DATA;
    output [31:0] PIPETX3DATA;
    output [31:0] PIPETX4DATA;
    output [31:0] PIPETX5DATA;
    output [31:0] PIPETX6DATA;
    output [31:0] PIPETX7DATA;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [3:0] CFGNEGOTIATEDWIDTH;
    output [3:0] CFGTPHSTTWRITEBYTEVALID;
    output [3:0] MICOMPLETIONRAMREADENABLEL;
    output [3:0] MICOMPLETIONRAMREADENABLEU;
    output [3:0] MICOMPLETIONRAMWRITEENABLEL;
    output [3:0] MICOMPLETIONRAMWRITEENABLEU;
    output [3:0] MIREQUESTRAMREADENABLE;
    output [3:0] MIREQUESTRAMWRITEENABLE;
    output [3:0] PCIERQSEQNUM;
    output [3:0] PIPERX0EQLPTXPRESET;
    output [3:0] PIPERX1EQLPTXPRESET;
    output [3:0] PIPERX2EQLPTXPRESET;
    output [3:0] PIPERX3EQLPTXPRESET;
    output [3:0] PIPERX4EQLPTXPRESET;
    output [3:0] PIPERX5EQLPTXPRESET;
    output [3:0] PIPERX6EQLPTXPRESET;
    output [3:0] PIPERX7EQLPTXPRESET;
    output [3:0] PIPETX0EQPRESET;
    output [3:0] PIPETX1EQPRESET;
    output [3:0] PIPETX2EQPRESET;
    output [3:0] PIPETX3EQPRESET;
    output [3:0] PIPETX4EQPRESET;
    output [3:0] PIPETX5EQPRESET;
    output [3:0] PIPETX6EQPRESET;
    output [3:0] PIPETX7EQPRESET;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output [4:0] CFGTPHSTTADDRESS;
    output [5:0] CFGFUNCTIONPOWERSTATE;
    output [5:0] CFGINTERRUPTMSIMMENABLE;
    output [5:0] CFGINTERRUPTMSIVFENABLE;
    output [5:0] CFGINTERRUPTMSIXVFENABLE;
    output [5:0] CFGINTERRUPTMSIXVFMASK;
    output [5:0] CFGLTSSMSTATE;
    output [5:0] CFGTPHSTMODE;
    output [5:0] CFGVFFLRINPROCESS;
    output [5:0] CFGVFTPHREQUESTERENABLE;
    output [5:0] PCIECQNPREQCOUNT;
    output [5:0] PCIERQTAG;
    output [5:0] PIPERX0EQLPLFFS;
    output [5:0] PIPERX1EQLPLFFS;
    output [5:0] PIPERX2EQLPLFFS;
    output [5:0] PIPERX3EQLPLFFS;
    output [5:0] PIPERX4EQLPLFFS;
    output [5:0] PIPERX5EQLPLFFS;
    output [5:0] PIPERX6EQLPLFFS;
    output [5:0] PIPERX7EQLPLFFS;
    output [5:0] PIPETX0EQDEEMPH;
    output [5:0] PIPETX1EQDEEMPH;
    output [5:0] PIPETX2EQDEEMPH;
    output [5:0] PIPETX3EQDEEMPH;
    output [5:0] PIPETX4EQDEEMPH;
    output [5:0] PIPETX5EQDEEMPH;
    output [5:0] PIPETX6EQDEEMPH;
    output [5:0] PIPETX7EQDEEMPH;
    output [71:0] MICOMPLETIONRAMWRITEDATAL;
    output [71:0] MICOMPLETIONRAMWRITEDATAU;
    output [74:0] MAXISRCTUSER;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output [7:0] CFGFCCPLH;
    output [7:0] CFGFCNPH;
    output [7:0] CFGFCPH;
    output [7:0] CFGFUNCTIONSTATUS;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [7:0] MAXISCQTKEEP;
    output [7:0] MAXISRCTKEEP;
    output [7:0] PLGEN3PCSRXSLIDE;
    output [84:0] MAXISCQTUSER;
    output [8:0] MIREPLAYRAMADDRESS;
    output [8:0] MIREQUESTRAMREADADDRESSA;
    output [8:0] MIREQUESTRAMREADADDRESSB;
    output [8:0] MIREQUESTRAMWRITEADDRESSA;
    output [8:0] MIREQUESTRAMWRITEADDRESSB;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [9:0] MICOMPLETIONRAMREADADDRESSAL;
    output [9:0] MICOMPLETIONRAMREADADDRESSAU;
    output [9:0] MICOMPLETIONRAMREADADDRESSBL;
    output [9:0] MICOMPLETIONRAMREADADDRESSBU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;
    input CFGCONFIGSPACEENABLE;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input CFGEXTREADDATAVALID;
    input CFGHOTRESETIN;
    input CFGINPUTUPDATEREQUEST;
    input CFGINTERRUPTMSITPHPRESENT;
    input CFGINTERRUPTMSIXINT;
    input CFGLINKTRAININGENABLE;
    input CFGMCUPDATEREQUEST;
    input CFGMGMTREAD;
    input CFGMGMTTYPE1CFGREGACCESS;
    input CFGMGMTWRITE;
    input CFGMSGTRANSMIT;
    input CFGPERFUNCTIONOUTPUTREQUEST;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input CFGTPHSTTREADDATAVALID;
    input CORECLK;
    input CORECLKMICOMPLETIONRAML;
    input CORECLKMICOMPLETIONRAMU;
    input CORECLKMIREPLAYRAM;
    input CORECLKMIREQUESTRAM;
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input PCIECQNPREQ;
    input PIPECLK;
    input PIPERESETN;
    input PIPERX0DATAVALID;
    input PIPERX0ELECIDLE;
    input PIPERX0EQDONE;
    input PIPERX0EQLPADAPTDONE;
    input PIPERX0EQLPLFFSSEL;
    input PIPERX0PHYSTATUS;
    input PIPERX0STARTBLOCK;
    input PIPERX0VALID;
    input PIPERX1DATAVALID;
    input PIPERX1ELECIDLE;
    input PIPERX1EQDONE;
    input PIPERX1EQLPADAPTDONE;
    input PIPERX1EQLPLFFSSEL;
    input PIPERX1PHYSTATUS;
    input PIPERX1STARTBLOCK;
    input PIPERX1VALID;
    input PIPERX2DATAVALID;
    input PIPERX2ELECIDLE;
    input PIPERX2EQDONE;
    input PIPERX2EQLPADAPTDONE;
    input PIPERX2EQLPLFFSSEL;
    input PIPERX2PHYSTATUS;
    input PIPERX2STARTBLOCK;
    input PIPERX2VALID;
    input PIPERX3DATAVALID;
    input PIPERX3ELECIDLE;
    input PIPERX3EQDONE;
    input PIPERX3EQLPADAPTDONE;
    input PIPERX3EQLPLFFSSEL;
    input PIPERX3PHYSTATUS;
    input PIPERX3STARTBLOCK;
    input PIPERX3VALID;
    input PIPERX4DATAVALID;
    input PIPERX4ELECIDLE;
    input PIPERX4EQDONE;
    input PIPERX4EQLPADAPTDONE;
    input PIPERX4EQLPLFFSSEL;
    input PIPERX4PHYSTATUS;
    input PIPERX4STARTBLOCK;
    input PIPERX4VALID;
    input PIPERX5DATAVALID;
    input PIPERX5ELECIDLE;
    input PIPERX5EQDONE;
    input PIPERX5EQLPADAPTDONE;
    input PIPERX5EQLPLFFSSEL;
    input PIPERX5PHYSTATUS;
    input PIPERX5STARTBLOCK;
    input PIPERX5VALID;
    input PIPERX6DATAVALID;
    input PIPERX6ELECIDLE;
    input PIPERX6EQDONE;
    input PIPERX6EQLPADAPTDONE;
    input PIPERX6EQLPLFFSSEL;
    input PIPERX6PHYSTATUS;
    input PIPERX6STARTBLOCK;
    input PIPERX6VALID;
    input PIPERX7DATAVALID;
    input PIPERX7ELECIDLE;
    input PIPERX7EQDONE;
    input PIPERX7EQLPADAPTDONE;
    input PIPERX7EQLPLFFSSEL;
    input PIPERX7PHYSTATUS;
    input PIPERX7STARTBLOCK;
    input PIPERX7VALID;
    input PIPETX0EQDONE;
    input PIPETX1EQDONE;
    input PIPETX2EQDONE;
    input PIPETX3EQDONE;
    input PIPETX4EQDONE;
    input PIPETX5EQDONE;
    input PIPETX6EQDONE;
    input PIPETX7EQDONE;
    input PLDISABLESCRAMBLER;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN3PCSDISABLE;
    input RECCLK;
    input RESETN;
    input SAXISCCTLAST;
    input SAXISCCTVALID;
    input SAXISRQTLAST;
    input SAXISRQTVALID;
    input USERCLK;
    input [10:0] DRPADDR;
    input [143:0] MICOMPLETIONRAMREADDATA;
    input [143:0] MIREPLAYRAMREADDATA;
    input [143:0] MIREQUESTRAMREADDATA;
    input [15:0] CFGDEVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [15:0] CFGVENDID;
    input [15:0] DRPDI;
    input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPETX0EQCOEFF;
    input [17:0] PIPETX1EQCOEFF;
    input [17:0] PIPETX2EQCOEFF;
    input [17:0] PIPETX3EQCOEFF;
    input [17:0] PIPETX4EQCOEFF;
    input [17:0] PIPETX5EQCOEFF;
    input [17:0] PIPETX6EQCOEFF;
    input [17:0] PIPETX7EQCOEFF;
    input [18:0] CFGMGMTADDR;
    input [1:0] CFGFLRDONE;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [1:0] CFGINTERRUPTPENDING;
    input [1:0] PIPERX0CHARISK;
    input [1:0] PIPERX0SYNCHEADER;
    input [1:0] PIPERX1CHARISK;
    input [1:0] PIPERX1SYNCHEADER;
    input [1:0] PIPERX2CHARISK;
    input [1:0] PIPERX2SYNCHEADER;
    input [1:0] PIPERX3CHARISK;
    input [1:0] PIPERX3SYNCHEADER;
    input [1:0] PIPERX4CHARISK;
    input [1:0] PIPERX4SYNCHEADER;
    input [1:0] PIPERX5CHARISK;
    input [1:0] PIPERX5SYNCHEADER;
    input [1:0] PIPERX6CHARISK;
    input [1:0] PIPERX6SYNCHEADER;
    input [1:0] PIPERX7CHARISK;
    input [1:0] PIPERX7SYNCHEADER;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input [255:0] SAXISCCTDATA;
    input [255:0] SAXISRQTDATA;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [2:0] CFGFCSEL;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [2:0] CFGPERFUNCSTATUSCONTROL;
    input [2:0] CFGPERFUNCTIONNUMBER;
    input [2:0] PIPERX0STATUS;
    input [2:0] PIPERX1STATUS;
    input [2:0] PIPERX2STATUS;
    input [2:0] PIPERX3STATUS;
    input [2:0] PIPERX4STATUS;
    input [2:0] PIPERX5STATUS;
    input [2:0] PIPERX6STATUS;
    input [2:0] PIPERX7STATUS;
    input [31:0] CFGEXTREADDATA;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input [31:0] CFGMGMTWRITEDATA;
    input [31:0] CFGMSGTRANSMITDATA;
    input [31:0] CFGTPHSTTREADDATA;
    input [31:0] PIPERX0DATA;
    input [31:0] PIPERX1DATA;
    input [31:0] PIPERX2DATA;
    input [31:0] PIPERX3DATA;
    input [31:0] PIPERX4DATA;
    input [31:0] PIPERX5DATA;
    input [31:0] PIPERX6DATA;
    input [31:0] PIPERX7DATA;
    input [32:0] SAXISCCTUSER;
    input [3:0] CFGINTERRUPTINT;
    input [3:0] CFGINTERRUPTMSISELECT;
    input [3:0] CFGMGMTBYTEENABLE;
    input [4:0] CFGDSDEVICENUMBER;
    input [59:0] SAXISRQTUSER;
    input [5:0] CFGVFFLRDONE;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input [63:0] CFGDSN;
    input [63:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [7:0] CFGDSBUSNUMBER;
    input [7:0] CFGDSPORTNUMBER;
    input [7:0] CFGREVID;
    input [7:0] PLGEN3PCSRXSYNCDONE;
    input [7:0] SAXISCCTKEEP;
    input [7:0] SAXISRQTKEEP;
    input [8:0] CFGINTERRUPTMSITPHSTTAG;
endmodule

module PCIE_3_1 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
    parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE = "FALSE";
    parameter DEBUG_PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF0_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_BIST_REGISTER = 8'h00;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter [15:0] PF0_DEVICE_ID = 16'h0000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF0_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
    parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF0_PB_CAP_VER = 4'h1;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter PF0_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF0_RBAR_NUM = 3'h1;
    parameter [7:0] PF0_REVISION_ID = 8'h00;
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF1_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_BIST_REGISTER = 8'h00;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [15:0] PF1_DEVICE_ID = 16'h0000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF1_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
    parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF1_PB_CAP_VER = 4'h1;
    parameter [7:0] PF1_PM_CAP_ID = 8'h01;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
    parameter PF1_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF1_RBAR_NUM = 3'h1;
    parameter [7:0] PF1_REVISION_ID = 8'h00;
    parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
    parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF1_TPHR_CAP_ENABLE = "FALSE";
    parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
    parameter PF2_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF2_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF2_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF2_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF2_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_BIST_REGISTER = 8'h00;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [15:0] PF2_DEVICE_ID = 16'h0000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF2_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF2_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF2_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF2_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF2_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF2_PB_CAP_NEXTPTR = 12'h000;
    parameter PF2_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF2_PB_CAP_VER = 4'h1;
    parameter [7:0] PF2_PM_CAP_ID = 8'h01;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF2_PM_CAP_VER_ID = 3'h3;
    parameter PF2_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF2_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF2_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF2_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF2_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF2_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF2_RBAR_NUM = 3'h1;
    parameter [7:0] PF2_REVISION_ID = 8'h00;
    parameter [4:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF2_SUBSYSTEM_ID = 16'h0000;
    parameter PF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF2_TPHR_CAP_ENABLE = "FALSE";
    parameter PF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF2_TPHR_CAP_VER = 4'h1;
    parameter PF3_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF3_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF3_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF3_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF3_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_BIST_REGISTER = 8'h00;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [15:0] PF3_DEVICE_ID = 16'h0000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF3_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF3_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF3_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF3_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF3_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF3_PB_CAP_NEXTPTR = 12'h000;
    parameter PF3_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF3_PB_CAP_VER = 4'h1;
    parameter [7:0] PF3_PM_CAP_ID = 8'h01;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF3_PM_CAP_VER_ID = 3'h3;
    parameter PF3_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF3_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF3_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF3_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF3_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF3_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF3_RBAR_NUM = 3'h1;
    parameter [7:0] PF3_REVISION_ID = 8'h00;
    parameter [4:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF3_SUBSYSTEM_ID = 16'h0000;
    parameter PF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF3_TPHR_CAP_ENABLE = "FALSE";
    parameter PF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF3_TPHR_CAP_VER = 4'h1;
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP = "TRUE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter PL_DISABLE_SCRAMBLING = "FALSE";
    parameter PL_DISABLE_SYNC_HEADER_FRAMING_ERROR = "FALSE";
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
    parameter [2:0] PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT = 3'h3;
    parameter [3:0] PL_EQ_DEFAULT_GEN3_TX_PRESET = 4'h4;
    parameter PL_EQ_PHASE01_RX_ADAPT = "FALSE";
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
    parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
    parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
    parameter integer PL_N_FTS_GEN1 = 255;
    parameter integer PL_N_FTS_GEN2 = 255;
    parameter integer PL_N_FTS_GEN3 = 255;
    parameter PL_REPORT_ALL_PHY_ERRORS = "TRUE";
    parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SRIOV_CAP_ENABLE = "FALSE";
    parameter TL_COMPLETION_RAM_SIZE_16K = "TRUE";
    parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [11:0] TL_CREDITS_CD = 12'h3E0;
    parameter [7:0] TL_CREDITS_CH = 8'h20;
    parameter [11:0] TL_CREDITS_NPD = 12'h028;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h198;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
    parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_MODE_ENABLE = "FALSE";
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TWO_LAYER_MODE_DLCMSM_ENABLE = "TRUE";
    parameter TWO_LAYER_MODE_ENABLE = "FALSE";
    parameter TWO_LAYER_MODE_WIDTH_256 = "TRUE";
    parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
    parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF0_PM_CAP_ID = 8'h01;
    parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
    parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF0_TPHR_CAP_ENABLE = "FALSE";
    parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF1_PM_CAP_ID = 8'h01;
    parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
    parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF1_TPHR_CAP_ENABLE = "FALSE";
    parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF2_PM_CAP_ID = 8'h01;
    parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
    parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF2_TPHR_CAP_ENABLE = "FALSE";
    parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF3_PM_CAP_ID = 8'h01;
    parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
    parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF3_TPHR_CAP_ENABLE = "FALSE";
    parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF4_PM_CAP_ID = 8'h01;
    parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
    parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF4_TPHR_CAP_ENABLE = "FALSE";
    parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF5_PM_CAP_ID = 8'h01;
    parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
    parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF5_TPHR_CAP_ENABLE = "FALSE";
    parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF6_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF6_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF6_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF6_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF6_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF6_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF6_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF6_PM_CAP_ID = 8'h01;
    parameter [7:0] VF6_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF6_PM_CAP_VER_ID = 3'h3;
    parameter VF6_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF6_TPHR_CAP_ENABLE = "FALSE";
    parameter VF6_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF6_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF6_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF6_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF6_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF6_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF7_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF7_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF7_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF7_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF7_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF7_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF7_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF7_PM_CAP_ID = 8'h01;
    parameter [7:0] VF7_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF7_PM_CAP_VER_ID = 3'h3;
    parameter VF7_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF7_TPHR_CAP_ENABLE = "FALSE";
    parameter VF7_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF7_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF7_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF7_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF7_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF7_TPHR_CAP_VER = 4'h1;
    output [2:0] CFGCURRENTSPEED;
    output [3:0] CFGDPASUBSTATECHANGE;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [7:0] CFGINTERRUPTMSIVFENABLE;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFAIL;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXSENT;
    output [7:0] CFGINTERRUPTMSIXVFENABLE;
    output [7:0] CFGINTERRUPTMSIXVFMASK;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output CFGLOCALERROR;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [2:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [3:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output [15:0] CFGPERFUNCSTATUSDATA;
    output CFGPERFUNCTIONUPDATEDONE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [3:0] CFGTPHFUNCTIONNUM;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [4:0] CFGTPHSTTADDRESS;
    output CFGTPHSTTREADENABLE;
    output [3:0] CFGTPHSTTWRITEBYTEVALID;
    output [31:0] CFGTPHSTTWRITEDATA;
    output CFGTPHSTTWRITEENABLE;
    output [7:0] CFGVFFLRINPROCESS;
    output [23:0] CFGVFPOWERSTATE;
    output [15:0] CFGVFSTATUS;
    output [7:0] CFGVFTPHREQUESTERENABLE;
    output [23:0] CFGVFTPHSTMODE;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [15:0] DBGDATAOUT;
    output DBGMCAPCSB;
    output [31:0] DBGMCAPDATA;
    output DBGMCAPEOS;
    output DBGMCAPERROR;
    output DBGMCAPMODE;
    output DBGMCAPRDATAVALID;
    output DBGMCAPRDWRB;
    output DBGMCAPRESET;
    output DBGPLDATABLOCKRECEIVEDAFTEREDS;
    output DBGPLGEN3FRAMINGERRORDETECTED;
    output DBGPLGEN3SYNCHEADERERRORDETECTED;
    output [7:0] DBGPLINFERREDRXELECTRICALIDLE;
    output [15:0] DRPDO;
    output DRPRDY;
    output LL2LMMASTERTLPSENT0;
    output LL2LMMASTERTLPSENT1;
    output [3:0] LL2LMMASTERTLPSENTTLPID0;
    output [3:0] LL2LMMASTERTLPSENTTLPID1;
    output [255:0] LL2LMMAXISRXTDATA;
    output [17:0] LL2LMMAXISRXTUSER;
    output [7:0] LL2LMMAXISRXTVALID;
    output [7:0] LL2LMSAXISTXTREADY;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [84:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [9:0] MICOMPLETIONRAMREADADDRESSAL;
    output [9:0] MICOMPLETIONRAMREADADDRESSAU;
    output [9:0] MICOMPLETIONRAMREADADDRESSBL;
    output [9:0] MICOMPLETIONRAMREADADDRESSBU;
    output [3:0] MICOMPLETIONRAMREADENABLEL;
    output [3:0] MICOMPLETIONRAMREADENABLEU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;
    output [71:0] MICOMPLETIONRAMWRITEDATAL;
    output [71:0] MICOMPLETIONRAMWRITEDATAU;
    output [3:0] MICOMPLETIONRAMWRITEENABLEL;
    output [3:0] MICOMPLETIONRAMWRITEENABLEU;
    output [8:0] MIREPLAYRAMADDRESS;
    output [1:0] MIREPLAYRAMREADENABLE;
    output [143:0] MIREPLAYRAMWRITEDATA;
    output [1:0] MIREPLAYRAMWRITEENABLE;
    output [8:0] MIREQUESTRAMREADADDRESSA;
    output [8:0] MIREQUESTRAMREADADDRESSB;
    output [3:0] MIREQUESTRAMREADENABLE;
    output [8:0] MIREQUESTRAMWRITEADDRESSA;
    output [8:0] MIREQUESTRAMWRITEADDRESSB;
    output [143:0] MIREQUESTRAMWRITEDATA;
    output [3:0] MIREQUESTRAMWRITEENABLE;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [3:0] PCIERQSEQNUM;
    output PCIERQSEQNUMVLD;
    output [5:0] PCIERQTAG;
    output [1:0] PCIERQTAGAV;
    output PCIERQTAGVLD;
    output [1:0] PCIETFCNPDAV;
    output [1:0] PCIETFCNPHAV;
    output [1:0] PIPERX0EQCONTROL;
    output [5:0] PIPERX0EQLPLFFS;
    output [3:0] PIPERX0EQLPTXPRESET;
    output [2:0] PIPERX0EQPRESET;
    output PIPERX0POLARITY;
    output [1:0] PIPERX1EQCONTROL;
    output [5:0] PIPERX1EQLPLFFS;
    output [3:0] PIPERX1EQLPTXPRESET;
    output [2:0] PIPERX1EQPRESET;
    output PIPERX1POLARITY;
    output [1:0] PIPERX2EQCONTROL;
    output [5:0] PIPERX2EQLPLFFS;
    output [3:0] PIPERX2EQLPTXPRESET;
    output [2:0] PIPERX2EQPRESET;
    output PIPERX2POLARITY;
    output [1:0] PIPERX3EQCONTROL;
    output [5:0] PIPERX3EQLPLFFS;
    output [3:0] PIPERX3EQLPTXPRESET;
    output [2:0] PIPERX3EQPRESET;
    output PIPERX3POLARITY;
    output [1:0] PIPERX4EQCONTROL;
    output [5:0] PIPERX4EQLPLFFS;
    output [3:0] PIPERX4EQLPTXPRESET;
    output [2:0] PIPERX4EQPRESET;
    output PIPERX4POLARITY;
    output [1:0] PIPERX5EQCONTROL;
    output [5:0] PIPERX5EQLPLFFS;
    output [3:0] PIPERX5EQLPTXPRESET;
    output [2:0] PIPERX5EQPRESET;
    output PIPERX5POLARITY;
    output [1:0] PIPERX6EQCONTROL;
    output [5:0] PIPERX6EQLPLFFS;
    output [3:0] PIPERX6EQLPTXPRESET;
    output [2:0] PIPERX6EQPRESET;
    output PIPERX6POLARITY;
    output [1:0] PIPERX7EQCONTROL;
    output [5:0] PIPERX7EQLPLFFS;
    output [3:0] PIPERX7EQLPTXPRESET;
    output [2:0] PIPERX7EQPRESET;
    output PIPERX7POLARITY;
    output [1:0] PIPETX0CHARISK;
    output PIPETX0COMPLIANCE;
    output [31:0] PIPETX0DATA;
    output PIPETX0DATAVALID;
    output PIPETX0DEEMPH;
    output PIPETX0ELECIDLE;
    output [1:0] PIPETX0EQCONTROL;
    output [5:0] PIPETX0EQDEEMPH;
    output [3:0] PIPETX0EQPRESET;
    output [2:0] PIPETX0MARGIN;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX0RATE;
    output PIPETX0RCVRDET;
    output PIPETX0RESET;
    output PIPETX0STARTBLOCK;
    output PIPETX0SWING;
    output [1:0] PIPETX0SYNCHEADER;
    output [1:0] PIPETX1CHARISK;
    output PIPETX1COMPLIANCE;
    output [31:0] PIPETX1DATA;
    output PIPETX1DATAVALID;
    output PIPETX1DEEMPH;
    output PIPETX1ELECIDLE;
    output [1:0] PIPETX1EQCONTROL;
    output [5:0] PIPETX1EQDEEMPH;
    output [3:0] PIPETX1EQPRESET;
    output [2:0] PIPETX1MARGIN;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX1RATE;
    output PIPETX1RCVRDET;
    output PIPETX1RESET;
    output PIPETX1STARTBLOCK;
    output PIPETX1SWING;
    output [1:0] PIPETX1SYNCHEADER;
    output [1:0] PIPETX2CHARISK;
    output PIPETX2COMPLIANCE;
    output [31:0] PIPETX2DATA;
    output PIPETX2DATAVALID;
    output PIPETX2DEEMPH;
    output PIPETX2ELECIDLE;
    output [1:0] PIPETX2EQCONTROL;
    output [5:0] PIPETX2EQDEEMPH;
    output [3:0] PIPETX2EQPRESET;
    output [2:0] PIPETX2MARGIN;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX2RATE;
    output PIPETX2RCVRDET;
    output PIPETX2RESET;
    output PIPETX2STARTBLOCK;
    output PIPETX2SWING;
    output [1:0] PIPETX2SYNCHEADER;
    output [1:0] PIPETX3CHARISK;
    output PIPETX3COMPLIANCE;
    output [31:0] PIPETX3DATA;
    output PIPETX3DATAVALID;
    output PIPETX3DEEMPH;
    output PIPETX3ELECIDLE;
    output [1:0] PIPETX3EQCONTROL;
    output [5:0] PIPETX3EQDEEMPH;
    output [3:0] PIPETX3EQPRESET;
    output [2:0] PIPETX3MARGIN;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX3RATE;
    output PIPETX3RCVRDET;
    output PIPETX3RESET;
    output PIPETX3STARTBLOCK;
    output PIPETX3SWING;
    output [1:0] PIPETX3SYNCHEADER;
    output [1:0] PIPETX4CHARISK;
    output PIPETX4COMPLIANCE;
    output [31:0] PIPETX4DATA;
    output PIPETX4DATAVALID;
    output PIPETX4DEEMPH;
    output PIPETX4ELECIDLE;
    output [1:0] PIPETX4EQCONTROL;
    output [5:0] PIPETX4EQDEEMPH;
    output [3:0] PIPETX4EQPRESET;
    output [2:0] PIPETX4MARGIN;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX4RATE;
    output PIPETX4RCVRDET;
    output PIPETX4RESET;
    output PIPETX4STARTBLOCK;
    output PIPETX4SWING;
    output [1:0] PIPETX4SYNCHEADER;
    output [1:0] PIPETX5CHARISK;
    output PIPETX5COMPLIANCE;
    output [31:0] PIPETX5DATA;
    output PIPETX5DATAVALID;
    output PIPETX5DEEMPH;
    output PIPETX5ELECIDLE;
    output [1:0] PIPETX5EQCONTROL;
    output [5:0] PIPETX5EQDEEMPH;
    output [3:0] PIPETX5EQPRESET;
    output [2:0] PIPETX5MARGIN;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX5RATE;
    output PIPETX5RCVRDET;
    output PIPETX5RESET;
    output PIPETX5STARTBLOCK;
    output PIPETX5SWING;
    output [1:0] PIPETX5SYNCHEADER;
    output [1:0] PIPETX6CHARISK;
    output PIPETX6COMPLIANCE;
    output [31:0] PIPETX6DATA;
    output PIPETX6DATAVALID;
    output PIPETX6DEEMPH;
    output PIPETX6ELECIDLE;
    output [1:0] PIPETX6EQCONTROL;
    output [5:0] PIPETX6EQDEEMPH;
    output [3:0] PIPETX6EQPRESET;
    output [2:0] PIPETX6MARGIN;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX6RATE;
    output PIPETX6RCVRDET;
    output PIPETX6RESET;
    output PIPETX6STARTBLOCK;
    output PIPETX6SWING;
    output [1:0] PIPETX6SYNCHEADER;
    output [1:0] PIPETX7CHARISK;
    output PIPETX7COMPLIANCE;
    output [31:0] PIPETX7DATA;
    output PIPETX7DATAVALID;
    output PIPETX7DEEMPH;
    output PIPETX7ELECIDLE;
    output [1:0] PIPETX7EQCONTROL;
    output [5:0] PIPETX7EQDEEMPH;
    output [3:0] PIPETX7EQPRESET;
    output [2:0] PIPETX7MARGIN;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PIPETX7RATE;
    output PIPETX7RCVRDET;
    output PIPETX7RESET;
    output PIPETX7STARTBLOCK;
    output PIPETX7SWING;
    output [1:0] PIPETX7SYNCHEADER;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [31:0] SPAREOUT;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVID;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [3:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [3:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [3:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [8:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [18:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTREAD;
    input CFGMGMTTYPE1CFGREGACCESS;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [2:0] CFGPERFUNCSTATUSCONTROL;
    input [3:0] CFGPERFUNCTIONNUMBER;
    input CFGPERFUNCTIONOUTPUTREQUEST;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [31:0] CFGTPHSTTREADDATA;
    input CFGTPHSTTREADDATAVALID;
    input [15:0] CFGVENDID;
    input [7:0] CFGVFFLRDONE;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKMICOMPLETIONRAML;
    input CORECLKMICOMPLETIONRAMU;
    input CORECLKMIREPLAYRAM;
    input CORECLKMIREQUESTRAM;
    input DBGCFGLOCALMGMTREGOVERRIDE;
    input [3:0] DBGDATASEL;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [13:0] LL2LMSAXISTXTUSER;
    input LL2LMSAXISTXTVALID;
    input [3:0] LL2LMTXTLPID0;
    input [3:0] LL2LMTXTLPID1;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [143:0] MICOMPLETIONRAMREADDATA;
    input [143:0] MIREPLAYRAMREADDATA;
    input [143:0] MIREQUESTRAMREADDATA;
    input PCIECQNPREQ;
    input PIPECLK;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX0CHARISK;
    input [31:0] PIPERX0DATA;
    input PIPERX0DATAVALID;
    input PIPERX0ELECIDLE;
    input PIPERX0EQDONE;
    input PIPERX0EQLPADAPTDONE;
    input PIPERX0EQLPLFFSSEL;
    input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
    input PIPERX0PHYSTATUS;
    input PIPERX0STARTBLOCK;
    input [2:0] PIPERX0STATUS;
    input [1:0] PIPERX0SYNCHEADER;
    input PIPERX0VALID;
    input [1:0] PIPERX1CHARISK;
    input [31:0] PIPERX1DATA;
    input PIPERX1DATAVALID;
    input PIPERX1ELECIDLE;
    input PIPERX1EQDONE;
    input PIPERX1EQLPADAPTDONE;
    input PIPERX1EQLPLFFSSEL;
    input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
    input PIPERX1PHYSTATUS;
    input PIPERX1STARTBLOCK;
    input [2:0] PIPERX1STATUS;
    input [1:0] PIPERX1SYNCHEADER;
    input PIPERX1VALID;
    input [1:0] PIPERX2CHARISK;
    input [31:0] PIPERX2DATA;
    input PIPERX2DATAVALID;
    input PIPERX2ELECIDLE;
    input PIPERX2EQDONE;
    input PIPERX2EQLPADAPTDONE;
    input PIPERX2EQLPLFFSSEL;
    input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
    input PIPERX2PHYSTATUS;
    input PIPERX2STARTBLOCK;
    input [2:0] PIPERX2STATUS;
    input [1:0] PIPERX2SYNCHEADER;
    input PIPERX2VALID;
    input [1:0] PIPERX3CHARISK;
    input [31:0] PIPERX3DATA;
    input PIPERX3DATAVALID;
    input PIPERX3ELECIDLE;
    input PIPERX3EQDONE;
    input PIPERX3EQLPADAPTDONE;
    input PIPERX3EQLPLFFSSEL;
    input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
    input PIPERX3PHYSTATUS;
    input PIPERX3STARTBLOCK;
    input [2:0] PIPERX3STATUS;
    input [1:0] PIPERX3SYNCHEADER;
    input PIPERX3VALID;
    input [1:0] PIPERX4CHARISK;
    input [31:0] PIPERX4DATA;
    input PIPERX4DATAVALID;
    input PIPERX4ELECIDLE;
    input PIPERX4EQDONE;
    input PIPERX4EQLPADAPTDONE;
    input PIPERX4EQLPLFFSSEL;
    input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
    input PIPERX4PHYSTATUS;
    input PIPERX4STARTBLOCK;
    input [2:0] PIPERX4STATUS;
    input [1:0] PIPERX4SYNCHEADER;
    input PIPERX4VALID;
    input [1:0] PIPERX5CHARISK;
    input [31:0] PIPERX5DATA;
    input PIPERX5DATAVALID;
    input PIPERX5ELECIDLE;
    input PIPERX5EQDONE;
    input PIPERX5EQLPADAPTDONE;
    input PIPERX5EQLPLFFSSEL;
    input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
    input PIPERX5PHYSTATUS;
    input PIPERX5STARTBLOCK;
    input [2:0] PIPERX5STATUS;
    input [1:0] PIPERX5SYNCHEADER;
    input PIPERX5VALID;
    input [1:0] PIPERX6CHARISK;
    input [31:0] PIPERX6DATA;
    input PIPERX6DATAVALID;
    input PIPERX6ELECIDLE;
    input PIPERX6EQDONE;
    input PIPERX6EQLPADAPTDONE;
    input PIPERX6EQLPLFFSSEL;
    input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
    input PIPERX6PHYSTATUS;
    input PIPERX6STARTBLOCK;
    input [2:0] PIPERX6STATUS;
    input [1:0] PIPERX6SYNCHEADER;
    input PIPERX6VALID;
    input [1:0] PIPERX7CHARISK;
    input [31:0] PIPERX7DATA;
    input PIPERX7DATAVALID;
    input PIPERX7ELECIDLE;
    input PIPERX7EQDONE;
    input PIPERX7EQLPADAPTDONE;
    input PIPERX7EQLPLFFSSEL;
    input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
    input PIPERX7PHYSTATUS;
    input PIPERX7STARTBLOCK;
    input [2:0] PIPERX7STATUS;
    input [1:0] PIPERX7SYNCHEADER;
    input PIPERX7VALID;
    input [17:0] PIPETX0EQCOEFF;
    input PIPETX0EQDONE;
    input [17:0] PIPETX1EQCOEFF;
    input PIPETX1EQDONE;
    input [17:0] PIPETX2EQCOEFF;
    input PIPETX2EQDONE;
    input [17:0] PIPETX3EQCOEFF;
    input PIPETX3EQDONE;
    input [17:0] PIPETX4EQCOEFF;
    input PIPETX4EQDONE;
    input [17:0] PIPETX5EQCOEFF;
    input PIPETX5EQDONE;
    input [17:0] PIPETX6EQCOEFF;
    input PIPETX6EQDONE;
    input [17:0] PIPETX7EQCOEFF;
    input PIPETX7EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input RESETN;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [59:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input [31:0] SPAREIN;
    input USERCLK;
endmodule

module PCIE40E4 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AUTO_FLR_RESPONSE = "FALSE";
    parameter [1:0] AXISTEN_IF_CC_ALIGNMENT_MODE = 2'h0;
    parameter [23:0] AXISTEN_IF_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] AXISTEN_IF_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [1:0] AXISTEN_IF_CQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_CQ_EN_POISONED_MEM_WR = "FALSE";
    parameter AXISTEN_IF_ENABLE_256_TAGS = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE = "FALSE";
    parameter AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK = "TRUE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_EXT_512 = "FALSE";
    parameter AXISTEN_IF_EXT_512_CC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_CQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_LEGACY_MODE_ENABLE = "FALSE";
    parameter AXISTEN_IF_MSIX_FROM_RAM_PIPELINE = "FALSE";
    parameter AXISTEN_IF_MSIX_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_MSIX_TO_RAM_PIPELINE = "FALSE";
    parameter [1:0] AXISTEN_IF_RC_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter [1:0] AXISTEN_IF_RQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT = "FALSE";
    parameter AXISTEN_IF_TX_PARITY_EN = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CFG_BYPASS_MODE_ENABLE = "FALSE";
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter [15:0] DEBUG_AXI4ST_SPARE = 16'h0000;
    parameter [7:0] DEBUG_AXIST_DISABLE_FEATURE_BIT = 8'h00;
    parameter [3:0] DEBUG_CAR_SPARE = 4'h0;
    parameter [15:0] DEBUG_CFG_SPARE = 16'h0000;
    parameter [15:0] DEBUG_LL_SPARE = 16'h0000;
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW = "FALSE";
    parameter DEBUG_PL_DISABLE_SCRAMBLING = "FALSE";
    parameter DEBUG_PL_SIM_RESET_LFSR = "FALSE";
    parameter [15:0] DEBUG_PL_SPARE = 16'h0000;
    parameter DEBUG_TL_DISABLE_FC_TIMEOUT = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [15:0] DEBUG_TL_SPARE = 16'h0000;
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter DSN_CAP_ENABLE = "FALSE";
    parameter EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter HEADER_TYPE_OVERRIDE = "FALSE";
    parameter IS_SWITCH_PORT = "FALSE";
    parameter LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter LL_DISABLE_SCHED_TX_NAK = "FALSE";
    parameter LL_REPLAY_FROM_RAM_PIPELINE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter LL_REPLAY_TO_RAM_PIPELINE = "FALSE";
    parameter LL_RX_TLP_PARITY_GEN = "TRUE";
    parameter LL_TX_TLP_PARITY_CHK = "TRUE";
    parameter [15:0] LL_USER_SPARE = 16'h0000;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h250;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4 = 7;
    parameter [0:0] PF0_LINK_CONTROL_RCB = 1'h0;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [5:0] PF0_MSIX_VECTOR_COUNT = 6'h04;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter PL_CFG_STATE_ROBUSTNESS_ENABLE = "TRUE";
    parameter PL_DEEMPH_SOURCE_SELECT = "TRUE";
    parameter PL_DESKEW_ON_SKIP_IN_GEN12 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_LANE_REVERSAL = "FALSE";
    parameter [1:0] PL_DISABLE_LFSR_UPDATE_ON_SKP = 2'h0;
    parameter PL_DISABLE_RETRAIN_ON_EB_ERROR = "FALSE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter [15:0] PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR = 16'h0000;
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter [1:0] PL_EQ_ADAPT_DISABLE_COEFF_CHECK = 2'h0;
    parameter [1:0] PL_EQ_ADAPT_DISABLE_PRESET_CHECK = 2'h0;
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter [1:0] PL_EQ_BYPASS_PHASE23 = 2'h0;
    parameter [5:0] PL_EQ_DEFAULT_RX_PRESET_HINT = 6'h33;
    parameter [7:0] PL_EQ_DEFAULT_TX_PRESET = 8'h44;
    parameter PL_EQ_DISABLE_MISMATCH_CHECK = "TRUE";
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE0 = 2'h0;
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE1 = 2'h0;
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter PL_EQ_TX_8G_EQ_TS2_ENABLE = "FALSE";
    parameter PL_EXIT_LOOPBACK_ON_EI_ENTRY = "TRUE";
    parameter PL_INFER_EI_DISABLE_LPBK_ACTIVE = "TRUE";
    parameter PL_INFER_EI_DISABLE_REC_RC = "FALSE";
    parameter PL_INFER_EI_DISABLE_REC_SPD = "FALSE";
    parameter [31:0] PL_LANE0_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE10_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE11_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE12_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE13_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE14_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE15_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE1_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE2_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE3_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE4_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE5_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE6_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE7_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE8_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE9_EQ_CONTROL = 32'h00003F00;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_SPEED = 4'h4;
    parameter [4:0] PL_LINK_CAP_MAX_LINK_WIDTH = 5'h08;
    parameter integer PL_N_FTS = 255;
    parameter PL_QUIESCE_GUARANTEE_DISABLE = "FALSE";
    parameter PL_REDO_EQ_SOURCE_SELECT = "TRUE";
    parameter [7:0] PL_REPORT_ALL_PHY_ERRORS = 8'h00;
    parameter [1:0] PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN4 = 4'h0;
    parameter [1:0] PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN4 = 4'h0;
    parameter [1:0] PL_RX_L0S_EXIT_TO_RECOVERY = 2'h0;
    parameter [1:0] PL_SIM_FAST_LINK_TRAINING = 2'h0;
    parameter PL_SRIS_ENABLE = "FALSE";
    parameter [6:0] PL_SRIS_SKPOS_GEN_SPD_VEC = 7'h00;
    parameter [6:0] PL_SRIS_SKPOS_REC_SPD_VEC = 7'h00;
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PL_USER_SPARE = 16'h0000;
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h1500;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h003E8;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000100;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h00000;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0100;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter SPARE_BIT0 = "FALSE";
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter SPARE_BIT3 = "FALSE";
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter [3:0] SRIOV_CAP_ENABLE = 4'h0;
    parameter TL2CFG_IF_PARITY_CHK = "TRUE";
    parameter [1:0] TL_COMPLETION_RAM_NUM_TLPS = 2'h0;
    parameter [1:0] TL_COMPLETION_RAM_SIZE = 2'h1;
    parameter [11:0] TL_CREDITS_CD = 12'h000;
    parameter [7:0] TL_CREDITS_CH = 8'h00;
    parameter [11:0] TL_CREDITS_NPD = 12'h004;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h0E0;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TIME = 5'h02;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT = 5'h08;
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter [0:0] TL_POSTED_RAM_SIZE = 1'h0;
    parameter TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TL_TX_TLP_STRADDLE_ENABLE = "FALSE";
    parameter TL_TX_TLP_TERMINATE_PARITY = "FALSE";
    parameter [15:0] TL_USER_SPARE = 16'h0000;
    parameter TPH_FROM_RAM_PIPELINE = "FALSE";
    parameter TPH_TO_RAM_PIPELINE = "FALSE";
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h80;
    parameter [11:0] VFG0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    output [7:0] AXIUSEROUT;
    output [7:0] CFGBUSNUMBER;
    output [1:0] CFGCURRENTSPEED;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXVECPENDINGSTATUS;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output [4:0] CFGLOCALERROROUT;
    output CFGLOCALERRORVALID;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [1:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [12:0] CFGMSIXRAMADDRESS;
    output CFGMSIXRAMREADENABLE;
    output [3:0] CFGMSIXRAMWRITEBYTEENABLE;
    output [35:0] CFGMSIXRAMWRITEDATA;
    output [2:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [1:0] CFGRXPMSTATE;
    output [11:0] CFGTPHRAMADDRESS;
    output CFGTPHRAMREADENABLE;
    output [3:0] CFGTPHRAMWRITEBYTEENABLE;
    output [35:0] CFGTPHRAMWRITEDATA;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [1:0] CFGTXPMSTATE;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [31:0] DBGCTRL0OUT;
    output [31:0] DBGCTRL1OUT;
    output [255:0] DBGDATA0OUT;
    output [255:0] DBGDATA1OUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [87:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [8:0] MIREPLAYRAMADDRESS0;
    output [8:0] MIREPLAYRAMADDRESS1;
    output MIREPLAYRAMREADENABLE0;
    output MIREPLAYRAMREADENABLE1;
    output [127:0] MIREPLAYRAMWRITEDATA0;
    output [127:0] MIREPLAYRAMWRITEDATA1;
    output MIREPLAYRAMWRITEENABLE0;
    output MIREPLAYRAMWRITEENABLE1;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS1;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE0;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE1;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS1;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA0;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA1;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE0;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS1;
    output MIRXPOSTEDREQUESTRAMREADENABLE0;
    output MIRXPOSTEDREQUESTRAMREADENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS1;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA0;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA1;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE0;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE1;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [5:0] PCIERQSEQNUM0;
    output [5:0] PCIERQSEQNUM1;
    output PCIERQSEQNUMVLD0;
    output PCIERQSEQNUMVLD1;
    output [7:0] PCIERQTAG0;
    output [7:0] PCIERQTAG1;
    output [3:0] PCIERQTAGAV;
    output PCIERQTAGVLD0;
    output PCIERQTAGVLD1;
    output [3:0] PCIETFCNPDAV;
    output [3:0] PCIETFCNPHAV;
    output [1:0] PIPERX00EQCONTROL;
    output PIPERX00POLARITY;
    output [1:0] PIPERX01EQCONTROL;
    output PIPERX01POLARITY;
    output [1:0] PIPERX02EQCONTROL;
    output PIPERX02POLARITY;
    output [1:0] PIPERX03EQCONTROL;
    output PIPERX03POLARITY;
    output [1:0] PIPERX04EQCONTROL;
    output PIPERX04POLARITY;
    output [1:0] PIPERX05EQCONTROL;
    output PIPERX05POLARITY;
    output [1:0] PIPERX06EQCONTROL;
    output PIPERX06POLARITY;
    output [1:0] PIPERX07EQCONTROL;
    output PIPERX07POLARITY;
    output [1:0] PIPERX08EQCONTROL;
    output PIPERX08POLARITY;
    output [1:0] PIPERX09EQCONTROL;
    output PIPERX09POLARITY;
    output [1:0] PIPERX10EQCONTROL;
    output PIPERX10POLARITY;
    output [1:0] PIPERX11EQCONTROL;
    output PIPERX11POLARITY;
    output [1:0] PIPERX12EQCONTROL;
    output PIPERX12POLARITY;
    output [1:0] PIPERX13EQCONTROL;
    output PIPERX13POLARITY;
    output [1:0] PIPERX14EQCONTROL;
    output PIPERX14POLARITY;
    output [1:0] PIPERX15EQCONTROL;
    output PIPERX15POLARITY;
    output [5:0] PIPERXEQLPLFFS;
    output [3:0] PIPERXEQLPTXPRESET;
    output [1:0] PIPETX00CHARISK;
    output PIPETX00COMPLIANCE;
    output [31:0] PIPETX00DATA;
    output PIPETX00DATAVALID;
    output PIPETX00ELECIDLE;
    output [1:0] PIPETX00EQCONTROL;
    output [5:0] PIPETX00EQDEEMPH;
    output [1:0] PIPETX00POWERDOWN;
    output PIPETX00STARTBLOCK;
    output [1:0] PIPETX00SYNCHEADER;
    output [1:0] PIPETX01CHARISK;
    output PIPETX01COMPLIANCE;
    output [31:0] PIPETX01DATA;
    output PIPETX01DATAVALID;
    output PIPETX01ELECIDLE;
    output [1:0] PIPETX01EQCONTROL;
    output [5:0] PIPETX01EQDEEMPH;
    output [1:0] PIPETX01POWERDOWN;
    output PIPETX01STARTBLOCK;
    output [1:0] PIPETX01SYNCHEADER;
    output [1:0] PIPETX02CHARISK;
    output PIPETX02COMPLIANCE;
    output [31:0] PIPETX02DATA;
    output PIPETX02DATAVALID;
    output PIPETX02ELECIDLE;
    output [1:0] PIPETX02EQCONTROL;
    output [5:0] PIPETX02EQDEEMPH;
    output [1:0] PIPETX02POWERDOWN;
    output PIPETX02STARTBLOCK;
    output [1:0] PIPETX02SYNCHEADER;
    output [1:0] PIPETX03CHARISK;
    output PIPETX03COMPLIANCE;
    output [31:0] PIPETX03DATA;
    output PIPETX03DATAVALID;
    output PIPETX03ELECIDLE;
    output [1:0] PIPETX03EQCONTROL;
    output [5:0] PIPETX03EQDEEMPH;
    output [1:0] PIPETX03POWERDOWN;
    output PIPETX03STARTBLOCK;
    output [1:0] PIPETX03SYNCHEADER;
    output [1:0] PIPETX04CHARISK;
    output PIPETX04COMPLIANCE;
    output [31:0] PIPETX04DATA;
    output PIPETX04DATAVALID;
    output PIPETX04ELECIDLE;
    output [1:0] PIPETX04EQCONTROL;
    output [5:0] PIPETX04EQDEEMPH;
    output [1:0] PIPETX04POWERDOWN;
    output PIPETX04STARTBLOCK;
    output [1:0] PIPETX04SYNCHEADER;
    output [1:0] PIPETX05CHARISK;
    output PIPETX05COMPLIANCE;
    output [31:0] PIPETX05DATA;
    output PIPETX05DATAVALID;
    output PIPETX05ELECIDLE;
    output [1:0] PIPETX05EQCONTROL;
    output [5:0] PIPETX05EQDEEMPH;
    output [1:0] PIPETX05POWERDOWN;
    output PIPETX05STARTBLOCK;
    output [1:0] PIPETX05SYNCHEADER;
    output [1:0] PIPETX06CHARISK;
    output PIPETX06COMPLIANCE;
    output [31:0] PIPETX06DATA;
    output PIPETX06DATAVALID;
    output PIPETX06ELECIDLE;
    output [1:0] PIPETX06EQCONTROL;
    output [5:0] PIPETX06EQDEEMPH;
    output [1:0] PIPETX06POWERDOWN;
    output PIPETX06STARTBLOCK;
    output [1:0] PIPETX06SYNCHEADER;
    output [1:0] PIPETX07CHARISK;
    output PIPETX07COMPLIANCE;
    output [31:0] PIPETX07DATA;
    output PIPETX07DATAVALID;
    output PIPETX07ELECIDLE;
    output [1:0] PIPETX07EQCONTROL;
    output [5:0] PIPETX07EQDEEMPH;
    output [1:0] PIPETX07POWERDOWN;
    output PIPETX07STARTBLOCK;
    output [1:0] PIPETX07SYNCHEADER;
    output [1:0] PIPETX08CHARISK;
    output PIPETX08COMPLIANCE;
    output [31:0] PIPETX08DATA;
    output PIPETX08DATAVALID;
    output PIPETX08ELECIDLE;
    output [1:0] PIPETX08EQCONTROL;
    output [5:0] PIPETX08EQDEEMPH;
    output [1:0] PIPETX08POWERDOWN;
    output PIPETX08STARTBLOCK;
    output [1:0] PIPETX08SYNCHEADER;
    output [1:0] PIPETX09CHARISK;
    output PIPETX09COMPLIANCE;
    output [31:0] PIPETX09DATA;
    output PIPETX09DATAVALID;
    output PIPETX09ELECIDLE;
    output [1:0] PIPETX09EQCONTROL;
    output [5:0] PIPETX09EQDEEMPH;
    output [1:0] PIPETX09POWERDOWN;
    output PIPETX09STARTBLOCK;
    output [1:0] PIPETX09SYNCHEADER;
    output [1:0] PIPETX10CHARISK;
    output PIPETX10COMPLIANCE;
    output [31:0] PIPETX10DATA;
    output PIPETX10DATAVALID;
    output PIPETX10ELECIDLE;
    output [1:0] PIPETX10EQCONTROL;
    output [5:0] PIPETX10EQDEEMPH;
    output [1:0] PIPETX10POWERDOWN;
    output PIPETX10STARTBLOCK;
    output [1:0] PIPETX10SYNCHEADER;
    output [1:0] PIPETX11CHARISK;
    output PIPETX11COMPLIANCE;
    output [31:0] PIPETX11DATA;
    output PIPETX11DATAVALID;
    output PIPETX11ELECIDLE;
    output [1:0] PIPETX11EQCONTROL;
    output [5:0] PIPETX11EQDEEMPH;
    output [1:0] PIPETX11POWERDOWN;
    output PIPETX11STARTBLOCK;
    output [1:0] PIPETX11SYNCHEADER;
    output [1:0] PIPETX12CHARISK;
    output PIPETX12COMPLIANCE;
    output [31:0] PIPETX12DATA;
    output PIPETX12DATAVALID;
    output PIPETX12ELECIDLE;
    output [1:0] PIPETX12EQCONTROL;
    output [5:0] PIPETX12EQDEEMPH;
    output [1:0] PIPETX12POWERDOWN;
    output PIPETX12STARTBLOCK;
    output [1:0] PIPETX12SYNCHEADER;
    output [1:0] PIPETX13CHARISK;
    output PIPETX13COMPLIANCE;
    output [31:0] PIPETX13DATA;
    output PIPETX13DATAVALID;
    output PIPETX13ELECIDLE;
    output [1:0] PIPETX13EQCONTROL;
    output [5:0] PIPETX13EQDEEMPH;
    output [1:0] PIPETX13POWERDOWN;
    output PIPETX13STARTBLOCK;
    output [1:0] PIPETX13SYNCHEADER;
    output [1:0] PIPETX14CHARISK;
    output PIPETX14COMPLIANCE;
    output [31:0] PIPETX14DATA;
    output PIPETX14DATAVALID;
    output PIPETX14ELECIDLE;
    output [1:0] PIPETX14EQCONTROL;
    output [5:0] PIPETX14EQDEEMPH;
    output [1:0] PIPETX14POWERDOWN;
    output PIPETX14STARTBLOCK;
    output [1:0] PIPETX14SYNCHEADER;
    output [1:0] PIPETX15CHARISK;
    output PIPETX15COMPLIANCE;
    output [31:0] PIPETX15DATA;
    output PIPETX15DATAVALID;
    output PIPETX15ELECIDLE;
    output [1:0] PIPETX15EQCONTROL;
    output [5:0] PIPETX15EQDEEMPH;
    output [1:0] PIPETX15POWERDOWN;
    output PIPETX15STARTBLOCK;
    output [1:0] PIPETX15SYNCHEADER;
    output PIPETXDEEMPH;
    output [2:0] PIPETXMARGIN;
    output [1:0] PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PIPETXSWING;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output PLGEN34EQMISMATCH;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [31:0] USERSPAREOUT;
    input [7:0] AXIUSERIN;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVIDPF0;
    input [15:0] CFGDEVIDPF1;
    input [15:0] CFGDEVIDPF2;
    input [15:0] CFGDEVIDPF3;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [7:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [1:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [1:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [7:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [1:0] CFGINTERRUPTMSIXVECPENDING;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [9:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTDEBUGACCESS;
    input [7:0] CFGMGMTFUNCTIONNUMBER;
    input CFGMGMTREAD;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [35:0] CFGMSIXRAMREADDATA;
    input CFGPMASPML1ENTRYREJECT;
    input CFGPMASPMTXL0SENTRYDISABLE;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVIDPF0;
    input [7:0] CFGREVIDPF1;
    input [7:0] CFGREVIDPF2;
    input [7:0] CFGREVIDPF3;
    input [15:0] CFGSUBSYSIDPF0;
    input [15:0] CFGSUBSYSIDPF1;
    input [15:0] CFGSUBSYSIDPF2;
    input [15:0] CFGSUBSYSIDPF3;
    input [15:0] CFGSUBSYSVENDID;
    input [35:0] CFGTPHRAMREADDATA;
    input [15:0] CFGVENDID;
    input CFGVFFLRDONE;
    input [7:0] CFGVFFLRFUNCNUM;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKMIREPLAYRAM0;
    input CORECLKMIREPLAYRAM1;
    input CORECLKMIRXCOMPLETIONRAM0;
    input CORECLKMIRXCOMPLETIONRAM1;
    input CORECLKMIRXPOSTEDREQUESTRAM0;
    input CORECLKMIRXPOSTEDREQUESTRAM1;
    input [5:0] DBGSEL0;
    input [5:0] DBGSEL1;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [5:0] MIREPLAYRAMERRCOR;
    input [5:0] MIREPLAYRAMERRUNCOR;
    input [127:0] MIREPLAYRAMREADDATA0;
    input [127:0] MIREPLAYRAMREADDATA1;
    input [11:0] MIRXCOMPLETIONRAMERRCOR;
    input [11:0] MIRXCOMPLETIONRAMERRUNCOR;
    input [143:0] MIRXCOMPLETIONRAMREADDATA0;
    input [143:0] MIRXCOMPLETIONRAMREADDATA1;
    input [5:0] MIRXPOSTEDREQUESTRAMERRCOR;
    input [5:0] MIRXPOSTEDREQUESTRAMERRUNCOR;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA0;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA1;
    input [1:0] PCIECOMPLDELIVERED;
    input [7:0] PCIECOMPLDELIVEREDTAG0;
    input [7:0] PCIECOMPLDELIVEREDTAG1;
    input [1:0] PCIECQNPREQ;
    input PCIECQNPUSERCREDITRCVD;
    input PCIECQPIPELINEEMPTY;
    input PCIEPOSTEDREQDELIVERED;
    input PIPECLK;
    input PIPECLKEN;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX00CHARISK;
    input [31:0] PIPERX00DATA;
    input PIPERX00DATAVALID;
    input PIPERX00ELECIDLE;
    input PIPERX00EQDONE;
    input PIPERX00EQLPADAPTDONE;
    input PIPERX00EQLPLFFSSEL;
    input [17:0] PIPERX00EQLPNEWTXCOEFFORPRESET;
    input PIPERX00PHYSTATUS;
    input [1:0] PIPERX00STARTBLOCK;
    input [2:0] PIPERX00STATUS;
    input [1:0] PIPERX00SYNCHEADER;
    input PIPERX00VALID;
    input [1:0] PIPERX01CHARISK;
    input [31:0] PIPERX01DATA;
    input PIPERX01DATAVALID;
    input PIPERX01ELECIDLE;
    input PIPERX01EQDONE;
    input PIPERX01EQLPADAPTDONE;
    input PIPERX01EQLPLFFSSEL;
    input [17:0] PIPERX01EQLPNEWTXCOEFFORPRESET;
    input PIPERX01PHYSTATUS;
    input [1:0] PIPERX01STARTBLOCK;
    input [2:0] PIPERX01STATUS;
    input [1:0] PIPERX01SYNCHEADER;
    input PIPERX01VALID;
    input [1:0] PIPERX02CHARISK;
    input [31:0] PIPERX02DATA;
    input PIPERX02DATAVALID;
    input PIPERX02ELECIDLE;
    input PIPERX02EQDONE;
    input PIPERX02EQLPADAPTDONE;
    input PIPERX02EQLPLFFSSEL;
    input [17:0] PIPERX02EQLPNEWTXCOEFFORPRESET;
    input PIPERX02PHYSTATUS;
    input [1:0] PIPERX02STARTBLOCK;
    input [2:0] PIPERX02STATUS;
    input [1:0] PIPERX02SYNCHEADER;
    input PIPERX02VALID;
    input [1:0] PIPERX03CHARISK;
    input [31:0] PIPERX03DATA;
    input PIPERX03DATAVALID;
    input PIPERX03ELECIDLE;
    input PIPERX03EQDONE;
    input PIPERX03EQLPADAPTDONE;
    input PIPERX03EQLPLFFSSEL;
    input [17:0] PIPERX03EQLPNEWTXCOEFFORPRESET;
    input PIPERX03PHYSTATUS;
    input [1:0] PIPERX03STARTBLOCK;
    input [2:0] PIPERX03STATUS;
    input [1:0] PIPERX03SYNCHEADER;
    input PIPERX03VALID;
    input [1:0] PIPERX04CHARISK;
    input [31:0] PIPERX04DATA;
    input PIPERX04DATAVALID;
    input PIPERX04ELECIDLE;
    input PIPERX04EQDONE;
    input PIPERX04EQLPADAPTDONE;
    input PIPERX04EQLPLFFSSEL;
    input [17:0] PIPERX04EQLPNEWTXCOEFFORPRESET;
    input PIPERX04PHYSTATUS;
    input [1:0] PIPERX04STARTBLOCK;
    input [2:0] PIPERX04STATUS;
    input [1:0] PIPERX04SYNCHEADER;
    input PIPERX04VALID;
    input [1:0] PIPERX05CHARISK;
    input [31:0] PIPERX05DATA;
    input PIPERX05DATAVALID;
    input PIPERX05ELECIDLE;
    input PIPERX05EQDONE;
    input PIPERX05EQLPADAPTDONE;
    input PIPERX05EQLPLFFSSEL;
    input [17:0] PIPERX05EQLPNEWTXCOEFFORPRESET;
    input PIPERX05PHYSTATUS;
    input [1:0] PIPERX05STARTBLOCK;
    input [2:0] PIPERX05STATUS;
    input [1:0] PIPERX05SYNCHEADER;
    input PIPERX05VALID;
    input [1:0] PIPERX06CHARISK;
    input [31:0] PIPERX06DATA;
    input PIPERX06DATAVALID;
    input PIPERX06ELECIDLE;
    input PIPERX06EQDONE;
    input PIPERX06EQLPADAPTDONE;
    input PIPERX06EQLPLFFSSEL;
    input [17:0] PIPERX06EQLPNEWTXCOEFFORPRESET;
    input PIPERX06PHYSTATUS;
    input [1:0] PIPERX06STARTBLOCK;
    input [2:0] PIPERX06STATUS;
    input [1:0] PIPERX06SYNCHEADER;
    input PIPERX06VALID;
    input [1:0] PIPERX07CHARISK;
    input [31:0] PIPERX07DATA;
    input PIPERX07DATAVALID;
    input PIPERX07ELECIDLE;
    input PIPERX07EQDONE;
    input PIPERX07EQLPADAPTDONE;
    input PIPERX07EQLPLFFSSEL;
    input [17:0] PIPERX07EQLPNEWTXCOEFFORPRESET;
    input PIPERX07PHYSTATUS;
    input [1:0] PIPERX07STARTBLOCK;
    input [2:0] PIPERX07STATUS;
    input [1:0] PIPERX07SYNCHEADER;
    input PIPERX07VALID;
    input [1:0] PIPERX08CHARISK;
    input [31:0] PIPERX08DATA;
    input PIPERX08DATAVALID;
    input PIPERX08ELECIDLE;
    input PIPERX08EQDONE;
    input PIPERX08EQLPADAPTDONE;
    input PIPERX08EQLPLFFSSEL;
    input [17:0] PIPERX08EQLPNEWTXCOEFFORPRESET;
    input PIPERX08PHYSTATUS;
    input [1:0] PIPERX08STARTBLOCK;
    input [2:0] PIPERX08STATUS;
    input [1:0] PIPERX08SYNCHEADER;
    input PIPERX08VALID;
    input [1:0] PIPERX09CHARISK;
    input [31:0] PIPERX09DATA;
    input PIPERX09DATAVALID;
    input PIPERX09ELECIDLE;
    input PIPERX09EQDONE;
    input PIPERX09EQLPADAPTDONE;
    input PIPERX09EQLPLFFSSEL;
    input [17:0] PIPERX09EQLPNEWTXCOEFFORPRESET;
    input PIPERX09PHYSTATUS;
    input [1:0] PIPERX09STARTBLOCK;
    input [2:0] PIPERX09STATUS;
    input [1:0] PIPERX09SYNCHEADER;
    input PIPERX09VALID;
    input [1:0] PIPERX10CHARISK;
    input [31:0] PIPERX10DATA;
    input PIPERX10DATAVALID;
    input PIPERX10ELECIDLE;
    input PIPERX10EQDONE;
    input PIPERX10EQLPADAPTDONE;
    input PIPERX10EQLPLFFSSEL;
    input [17:0] PIPERX10EQLPNEWTXCOEFFORPRESET;
    input PIPERX10PHYSTATUS;
    input [1:0] PIPERX10STARTBLOCK;
    input [2:0] PIPERX10STATUS;
    input [1:0] PIPERX10SYNCHEADER;
    input PIPERX10VALID;
    input [1:0] PIPERX11CHARISK;
    input [31:0] PIPERX11DATA;
    input PIPERX11DATAVALID;
    input PIPERX11ELECIDLE;
    input PIPERX11EQDONE;
    input PIPERX11EQLPADAPTDONE;
    input PIPERX11EQLPLFFSSEL;
    input [17:0] PIPERX11EQLPNEWTXCOEFFORPRESET;
    input PIPERX11PHYSTATUS;
    input [1:0] PIPERX11STARTBLOCK;
    input [2:0] PIPERX11STATUS;
    input [1:0] PIPERX11SYNCHEADER;
    input PIPERX11VALID;
    input [1:0] PIPERX12CHARISK;
    input [31:0] PIPERX12DATA;
    input PIPERX12DATAVALID;
    input PIPERX12ELECIDLE;
    input PIPERX12EQDONE;
    input PIPERX12EQLPADAPTDONE;
    input PIPERX12EQLPLFFSSEL;
    input [17:0] PIPERX12EQLPNEWTXCOEFFORPRESET;
    input PIPERX12PHYSTATUS;
    input [1:0] PIPERX12STARTBLOCK;
    input [2:0] PIPERX12STATUS;
    input [1:0] PIPERX12SYNCHEADER;
    input PIPERX12VALID;
    input [1:0] PIPERX13CHARISK;
    input [31:0] PIPERX13DATA;
    input PIPERX13DATAVALID;
    input PIPERX13ELECIDLE;
    input PIPERX13EQDONE;
    input PIPERX13EQLPADAPTDONE;
    input PIPERX13EQLPLFFSSEL;
    input [17:0] PIPERX13EQLPNEWTXCOEFFORPRESET;
    input PIPERX13PHYSTATUS;
    input [1:0] PIPERX13STARTBLOCK;
    input [2:0] PIPERX13STATUS;
    input [1:0] PIPERX13SYNCHEADER;
    input PIPERX13VALID;
    input [1:0] PIPERX14CHARISK;
    input [31:0] PIPERX14DATA;
    input PIPERX14DATAVALID;
    input PIPERX14ELECIDLE;
    input PIPERX14EQDONE;
    input PIPERX14EQLPADAPTDONE;
    input PIPERX14EQLPLFFSSEL;
    input [17:0] PIPERX14EQLPNEWTXCOEFFORPRESET;
    input PIPERX14PHYSTATUS;
    input [1:0] PIPERX14STARTBLOCK;
    input [2:0] PIPERX14STATUS;
    input [1:0] PIPERX14SYNCHEADER;
    input PIPERX14VALID;
    input [1:0] PIPERX15CHARISK;
    input [31:0] PIPERX15DATA;
    input PIPERX15DATAVALID;
    input PIPERX15ELECIDLE;
    input PIPERX15EQDONE;
    input PIPERX15EQLPADAPTDONE;
    input PIPERX15EQLPLFFSSEL;
    input [17:0] PIPERX15EQLPNEWTXCOEFFORPRESET;
    input PIPERX15PHYSTATUS;
    input [1:0] PIPERX15STARTBLOCK;
    input [2:0] PIPERX15STATUS;
    input [1:0] PIPERX15SYNCHEADER;
    input PIPERX15VALID;
    input [17:0] PIPETX00EQCOEFF;
    input PIPETX00EQDONE;
    input [17:0] PIPETX01EQCOEFF;
    input PIPETX01EQDONE;
    input [17:0] PIPETX02EQCOEFF;
    input PIPETX02EQDONE;
    input [17:0] PIPETX03EQCOEFF;
    input PIPETX03EQDONE;
    input [17:0] PIPETX04EQCOEFF;
    input PIPETX04EQDONE;
    input [17:0] PIPETX05EQCOEFF;
    input PIPETX05EQDONE;
    input [17:0] PIPETX06EQCOEFF;
    input PIPETX06EQDONE;
    input [17:0] PIPETX07EQCOEFF;
    input PIPETX07EQDONE;
    input [17:0] PIPETX08EQCOEFF;
    input PIPETX08EQDONE;
    input [17:0] PIPETX09EQCOEFF;
    input PIPETX09EQDONE;
    input [17:0] PIPETX10EQCOEFF;
    input PIPETX10EQDONE;
    input [17:0] PIPETX11EQCOEFF;
    input PIPETX11EQDONE;
    input [17:0] PIPETX12EQCOEFF;
    input PIPETX12EQDONE;
    input [17:0] PIPETX13EQCOEFF;
    input PIPETX13EQDONE;
    input [17:0] PIPETX14EQCOEFF;
    input PIPETX14EQDONE;
    input [17:0] PIPETX15EQCOEFF;
    input PIPETX15EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input PLGEN34REDOEQSPEED;
    input PLGEN34REDOEQUALIZATION;
    input RESETN;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [61:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input USERCLK;
    input USERCLK2;
    input USERCLKEN;
    input [31:0] USERSPAREIN;
endmodule

module EMAC (...);
    parameter EMAC0_MODE = "RGMII";
    parameter EMAC1_MODE = "RGMII";
    output DCRHOSTDONEIR;
    output EMAC0CLIENTANINTERRUPT;
    output EMAC0CLIENTRXBADFRAME;
    output EMAC0CLIENTRXCLIENTCLKOUT;
    output EMAC0CLIENTRXDVLD;
    output EMAC0CLIENTRXDVLDMSW;
    output EMAC0CLIENTRXDVREG6;
    output EMAC0CLIENTRXFRAMEDROP;
    output EMAC0CLIENTRXGOODFRAME;
    output EMAC0CLIENTRXSTATSBYTEVLD;
    output EMAC0CLIENTRXSTATSVLD;
    output EMAC0CLIENTTXACK;
    output EMAC0CLIENTTXCLIENTCLKOUT;
    output EMAC0CLIENTTXCOLLISION;
    output EMAC0CLIENTTXGMIIMIICLKOUT;
    output EMAC0CLIENTTXRETRANSMIT;
    output EMAC0CLIENTTXSTATS;
    output EMAC0CLIENTTXSTATSBYTEVLD;
    output EMAC0CLIENTTXSTATSVLD;
    output EMAC0PHYENCOMMAALIGN;
    output EMAC0PHYLOOPBACKMSB;
    output EMAC0PHYMCLKOUT;
    output EMAC0PHYMDOUT;
    output EMAC0PHYMDTRI;
    output EMAC0PHYMGTRXRESET;
    output EMAC0PHYMGTTXRESET;
    output EMAC0PHYPOWERDOWN;
    output EMAC0PHYSYNCACQSTATUS;
    output EMAC0PHYTXCHARDISPMODE;
    output EMAC0PHYTXCHARDISPVAL;
    output EMAC0PHYTXCHARISK;
    output EMAC0PHYTXCLK;
    output EMAC0PHYTXEN;
    output EMAC0PHYTXER;
    output EMAC1CLIENTANINTERRUPT;
    output EMAC1CLIENTRXBADFRAME;
    output EMAC1CLIENTRXCLIENTCLKOUT;
    output EMAC1CLIENTRXDVLD;
    output EMAC1CLIENTRXDVLDMSW;
    output EMAC1CLIENTRXDVREG6;
    output EMAC1CLIENTRXFRAMEDROP;
    output EMAC1CLIENTRXGOODFRAME;
    output EMAC1CLIENTRXSTATSBYTEVLD;
    output EMAC1CLIENTRXSTATSVLD;
    output EMAC1CLIENTTXACK;
    output EMAC1CLIENTTXCLIENTCLKOUT;
    output EMAC1CLIENTTXCOLLISION;
    output EMAC1CLIENTTXGMIIMIICLKOUT;
    output EMAC1CLIENTTXRETRANSMIT;
    output EMAC1CLIENTTXSTATS;
    output EMAC1CLIENTTXSTATSBYTEVLD;
    output EMAC1CLIENTTXSTATSVLD;
    output EMAC1PHYENCOMMAALIGN;
    output EMAC1PHYLOOPBACKMSB;
    output EMAC1PHYMCLKOUT;
    output EMAC1PHYMDOUT;
    output EMAC1PHYMDTRI;
    output EMAC1PHYMGTRXRESET;
    output EMAC1PHYMGTTXRESET;
    output EMAC1PHYPOWERDOWN;
    output EMAC1PHYSYNCACQSTATUS;
    output EMAC1PHYTXCHARDISPMODE;
    output EMAC1PHYTXCHARDISPVAL;
    output EMAC1PHYTXCHARISK;
    output EMAC1PHYTXCLK;
    output EMAC1PHYTXEN;
    output EMAC1PHYTXER;
    output EMACDCRACK;
    output HOSTMIIMRDY;
    output [0:31] EMACDCRDBUS;
    output [15:0] EMAC0CLIENTRXD;
    output [15:0] EMAC1CLIENTRXD;
    output [31:0] HOSTRDDATA;
    output [6:0] EMAC0CLIENTRXSTATS;
    output [6:0] EMAC1CLIENTRXSTATS;
    output [7:0] EMAC0PHYTXD;
    output [7:0] EMAC1PHYTXD;
    input CLIENTEMAC0DCMLOCKED;
    input CLIENTEMAC0PAUSEREQ;
    input CLIENTEMAC0RXCLIENTCLKIN;
    input CLIENTEMAC0TXCLIENTCLKIN;
    input CLIENTEMAC0TXDVLD;
    input CLIENTEMAC0TXDVLDMSW;
    input CLIENTEMAC0TXFIRSTBYTE;
    input CLIENTEMAC0TXGMIIMIICLKIN;
    input CLIENTEMAC0TXUNDERRUN;
    input CLIENTEMAC1DCMLOCKED;
    input CLIENTEMAC1PAUSEREQ;
    input CLIENTEMAC1RXCLIENTCLKIN;
    input CLIENTEMAC1TXCLIENTCLKIN;
    input CLIENTEMAC1TXDVLD;
    input CLIENTEMAC1TXDVLDMSW;
    input CLIENTEMAC1TXFIRSTBYTE;
    input CLIENTEMAC1TXGMIIMIICLKIN;
    input CLIENTEMAC1TXUNDERRUN;
    input DCREMACCLK;
    input DCREMACENABLE;
    input DCREMACREAD;
    input DCREMACWRITE;
    input HOSTCLK;
    input HOSTEMAC1SEL;
    input HOSTMIIMSEL;
    input HOSTREQ;
    input PHYEMAC0COL;
    input PHYEMAC0CRS;
    input PHYEMAC0GTXCLK;
    input PHYEMAC0MCLKIN;
    input PHYEMAC0MDIN;
    input PHYEMAC0MIITXCLK;
    input PHYEMAC0RXBUFERR;
    input PHYEMAC0RXCHARISCOMMA;
    input PHYEMAC0RXCHARISK;
    input PHYEMAC0RXCHECKINGCRC;
    input PHYEMAC0RXCLK;
    input PHYEMAC0RXCOMMADET;
    input PHYEMAC0RXDISPERR;
    input PHYEMAC0RXDV;
    input PHYEMAC0RXER;
    input PHYEMAC0RXNOTINTABLE;
    input PHYEMAC0RXRUNDISP;
    input PHYEMAC0SIGNALDET;
    input PHYEMAC0TXBUFERR;
    input PHYEMAC1COL;
    input PHYEMAC1CRS;
    input PHYEMAC1GTXCLK;
    input PHYEMAC1MCLKIN;
    input PHYEMAC1MDIN;
    input PHYEMAC1MIITXCLK;
    input PHYEMAC1RXBUFERR;
    input PHYEMAC1RXCHARISCOMMA;
    input PHYEMAC1RXCHARISK;
    input PHYEMAC1RXCHECKINGCRC;
    input PHYEMAC1RXCLK;
    input PHYEMAC1RXCOMMADET;
    input PHYEMAC1RXDISPERR;
    input PHYEMAC1RXDV;
    input PHYEMAC1RXER;
    input PHYEMAC1RXNOTINTABLE;
    input PHYEMAC1RXRUNDISP;
    input PHYEMAC1SIGNALDET;
    input PHYEMAC1TXBUFERR;
    input RESET;
    input [0:31] DCREMACDBUS;
    input [15:0] CLIENTEMAC0PAUSEVAL;
    input [15:0] CLIENTEMAC0TXD;
    input [15:0] CLIENTEMAC1PAUSEVAL;
    input [15:0] CLIENTEMAC1TXD;
    input [1:0] HOSTOPCODE;
    input [1:0] PHYEMAC0RXBUFSTATUS;
    input [1:0] PHYEMAC0RXLOSSOFSYNC;
    input [1:0] PHYEMAC1RXBUFSTATUS;
    input [1:0] PHYEMAC1RXLOSSOFSYNC;
    input [2:0] PHYEMAC0RXCLKCORCNT;
    input [2:0] PHYEMAC1RXCLKCORCNT;
    input [31:0] HOSTWRDATA;
    input [47:0] TIEEMAC0UNICASTADDR;
    input [47:0] TIEEMAC1UNICASTADDR;
    input [4:0] PHYEMAC0PHYAD;
    input [4:0] PHYEMAC1PHYAD;
    input [79:0] TIEEMAC0CONFIGVEC;
    input [79:0] TIEEMAC1CONFIGVEC;
    input [7:0] CLIENTEMAC0TXIFGDELAY;
    input [7:0] CLIENTEMAC1TXIFGDELAY;
    input [7:0] PHYEMAC0RXD;
    input [7:0] PHYEMAC1RXD;
    input [8:9] DCREMACABUS;
    input [9:0] HOSTADDR;
endmodule

module TEMAC (...);
    parameter EMAC0_1000BASEX_ENABLE = "FALSE";
    parameter EMAC0_ADDRFILTER_ENABLE = "FALSE";
    parameter EMAC0_BYTEPHY = "FALSE";
    parameter EMAC0_CONFIGVEC_79 = "FALSE";
    parameter EMAC0_GTLOOPBACK = "FALSE";
    parameter EMAC0_HOST_ENABLE = "FALSE";
    parameter EMAC0_LTCHECK_DISABLE = "FALSE";
    parameter EMAC0_MDIO_ENABLE = "FALSE";
    parameter EMAC0_PHYINITAUTONEG_ENABLE = "FALSE";
    parameter EMAC0_PHYISOLATE = "FALSE";
    parameter EMAC0_PHYLOOPBACKMSB = "FALSE";
    parameter EMAC0_PHYPOWERDOWN = "FALSE";
    parameter EMAC0_PHYRESET = "FALSE";
    parameter EMAC0_RGMII_ENABLE = "FALSE";
    parameter EMAC0_RX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC0_RXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC0_RXHALFDUPLEX = "FALSE";
    parameter EMAC0_RXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC0_RXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC0_RXRESET = "FALSE";
    parameter EMAC0_RXVLAN_ENABLE = "FALSE";
    parameter EMAC0_RX_ENABLE = "FALSE";
    parameter EMAC0_SGMII_ENABLE = "FALSE";
    parameter EMAC0_SPEED_LSB = "FALSE";
    parameter EMAC0_SPEED_MSB = "FALSE";
    parameter EMAC0_TX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC0_TXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC0_TXHALFDUPLEX = "FALSE";
    parameter EMAC0_TXIFGADJUST_ENABLE = "FALSE";
    parameter EMAC0_TXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC0_TXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC0_TXRESET = "FALSE";
    parameter EMAC0_TXVLAN_ENABLE = "FALSE";
    parameter EMAC0_TX_ENABLE = "FALSE";
    parameter EMAC0_UNIDIRECTION_ENABLE = "FALSE";
    parameter EMAC0_USECLKEN = "FALSE";
    parameter EMAC1_1000BASEX_ENABLE = "FALSE";
    parameter EMAC1_ADDRFILTER_ENABLE = "FALSE";
    parameter EMAC1_BYTEPHY = "FALSE";
    parameter EMAC1_CONFIGVEC_79 = "FALSE";
    parameter EMAC1_GTLOOPBACK = "FALSE";
    parameter EMAC1_HOST_ENABLE = "FALSE";
    parameter EMAC1_LTCHECK_DISABLE = "FALSE";
    parameter EMAC1_MDIO_ENABLE = "FALSE";
    parameter EMAC1_PHYINITAUTONEG_ENABLE = "FALSE";
    parameter EMAC1_PHYISOLATE = "FALSE";
    parameter EMAC1_PHYLOOPBACKMSB = "FALSE";
    parameter EMAC1_PHYPOWERDOWN = "FALSE";
    parameter EMAC1_PHYRESET = "FALSE";
    parameter EMAC1_RGMII_ENABLE = "FALSE";
    parameter EMAC1_RX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC1_RXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC1_RXHALFDUPLEX = "FALSE";
    parameter EMAC1_RXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC1_RXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC1_RXRESET = "FALSE";
    parameter EMAC1_RXVLAN_ENABLE = "FALSE";
    parameter EMAC1_RX_ENABLE = "FALSE";
    parameter EMAC1_SGMII_ENABLE = "FALSE";
    parameter EMAC1_SPEED_LSB = "FALSE";
    parameter EMAC1_SPEED_MSB = "FALSE";
    parameter EMAC1_TX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC1_TXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC1_TXHALFDUPLEX = "FALSE";
    parameter EMAC1_TXIFGADJUST_ENABLE = "FALSE";
    parameter EMAC1_TXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC1_TXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC1_TXRESET = "FALSE";
    parameter EMAC1_TXVLAN_ENABLE = "FALSE";
    parameter EMAC1_TX_ENABLE = "FALSE";
    parameter EMAC1_UNIDIRECTION_ENABLE = "FALSE";
    parameter EMAC1_USECLKEN = "FALSE";
    parameter [0:7] EMAC0_DCRBASEADDR = 8'h00;
    parameter [0:7] EMAC1_DCRBASEADDR = 8'h00;
    parameter [47:0] EMAC0_PAUSEADDR = 48'h000000000000;
    parameter [47:0] EMAC0_UNICASTADDR = 48'h000000000000;
    parameter [47:0] EMAC1_PAUSEADDR = 48'h000000000000;
    parameter [47:0] EMAC1_UNICASTADDR = 48'h000000000000;
    parameter [8:0] EMAC0_LINKTIMERVAL = 9'h000;
    parameter [8:0] EMAC1_LINKTIMERVAL = 9'h000;
    output DCRHOSTDONEIR;
    output EMAC0CLIENTANINTERRUPT;
    output EMAC0CLIENTRXBADFRAME;
    output EMAC0CLIENTRXCLIENTCLKOUT;
    output EMAC0CLIENTRXDVLD;
    output EMAC0CLIENTRXDVLDMSW;
    output EMAC0CLIENTRXFRAMEDROP;
    output EMAC0CLIENTRXGOODFRAME;
    output EMAC0CLIENTRXSTATSBYTEVLD;
    output EMAC0CLIENTRXSTATSVLD;
    output EMAC0CLIENTTXACK;
    output EMAC0CLIENTTXCLIENTCLKOUT;
    output EMAC0CLIENTTXCOLLISION;
    output EMAC0CLIENTTXRETRANSMIT;
    output EMAC0CLIENTTXSTATS;
    output EMAC0CLIENTTXSTATSBYTEVLD;
    output EMAC0CLIENTTXSTATSVLD;
    output EMAC0PHYENCOMMAALIGN;
    output EMAC0PHYLOOPBACKMSB;
    output EMAC0PHYMCLKOUT;
    output EMAC0PHYMDOUT;
    output EMAC0PHYMDTRI;
    output EMAC0PHYMGTRXRESET;
    output EMAC0PHYMGTTXRESET;
    output EMAC0PHYPOWERDOWN;
    output EMAC0PHYSYNCACQSTATUS;
    output EMAC0PHYTXCHARDISPMODE;
    output EMAC0PHYTXCHARDISPVAL;
    output EMAC0PHYTXCHARISK;
    output EMAC0PHYTXCLK;
    output EMAC0PHYTXEN;
    output EMAC0PHYTXER;
    output EMAC0PHYTXGMIIMIICLKOUT;
    output EMAC0SPEEDIS10100;
    output EMAC1CLIENTANINTERRUPT;
    output EMAC1CLIENTRXBADFRAME;
    output EMAC1CLIENTRXCLIENTCLKOUT;
    output EMAC1CLIENTRXDVLD;
    output EMAC1CLIENTRXDVLDMSW;
    output EMAC1CLIENTRXFRAMEDROP;
    output EMAC1CLIENTRXGOODFRAME;
    output EMAC1CLIENTRXSTATSBYTEVLD;
    output EMAC1CLIENTRXSTATSVLD;
    output EMAC1CLIENTTXACK;
    output EMAC1CLIENTTXCLIENTCLKOUT;
    output EMAC1CLIENTTXCOLLISION;
    output EMAC1CLIENTTXRETRANSMIT;
    output EMAC1CLIENTTXSTATS;
    output EMAC1CLIENTTXSTATSBYTEVLD;
    output EMAC1CLIENTTXSTATSVLD;
    output EMAC1PHYENCOMMAALIGN;
    output EMAC1PHYLOOPBACKMSB;
    output EMAC1PHYMCLKOUT;
    output EMAC1PHYMDOUT;
    output EMAC1PHYMDTRI;
    output EMAC1PHYMGTRXRESET;
    output EMAC1PHYMGTTXRESET;
    output EMAC1PHYPOWERDOWN;
    output EMAC1PHYSYNCACQSTATUS;
    output EMAC1PHYTXCHARDISPMODE;
    output EMAC1PHYTXCHARDISPVAL;
    output EMAC1PHYTXCHARISK;
    output EMAC1PHYTXCLK;
    output EMAC1PHYTXEN;
    output EMAC1PHYTXER;
    output EMAC1PHYTXGMIIMIICLKOUT;
    output EMAC1SPEEDIS10100;
    output EMACDCRACK;
    output HOSTMIIMRDY;
    output [0:31] EMACDCRDBUS;
    output [15:0] EMAC0CLIENTRXD;
    output [15:0] EMAC1CLIENTRXD;
    output [31:0] HOSTRDDATA;
    output [6:0] EMAC0CLIENTRXSTATS;
    output [6:0] EMAC1CLIENTRXSTATS;
    output [7:0] EMAC0PHYTXD;
    output [7:0] EMAC1PHYTXD;
    input CLIENTEMAC0DCMLOCKED;
    input CLIENTEMAC0PAUSEREQ;
    input CLIENTEMAC0RXCLIENTCLKIN;
    input CLIENTEMAC0TXCLIENTCLKIN;
    input CLIENTEMAC0TXDVLD;
    input CLIENTEMAC0TXDVLDMSW;
    input CLIENTEMAC0TXFIRSTBYTE;
    input CLIENTEMAC0TXUNDERRUN;
    input CLIENTEMAC1DCMLOCKED;
    input CLIENTEMAC1PAUSEREQ;
    input CLIENTEMAC1RXCLIENTCLKIN;
    input CLIENTEMAC1TXCLIENTCLKIN;
    input CLIENTEMAC1TXDVLD;
    input CLIENTEMAC1TXDVLDMSW;
    input CLIENTEMAC1TXFIRSTBYTE;
    input CLIENTEMAC1TXUNDERRUN;
    input DCREMACCLK;
    input DCREMACENABLE;
    input DCREMACREAD;
    input DCREMACWRITE;
    input HOSTCLK;
    input HOSTEMAC1SEL;
    input HOSTMIIMSEL;
    input HOSTREQ;
    input PHYEMAC0COL;
    input PHYEMAC0CRS;
    input PHYEMAC0GTXCLK;
    input PHYEMAC0MCLKIN;
    input PHYEMAC0MDIN;
    input PHYEMAC0MIITXCLK;
    input PHYEMAC0RXBUFERR;
    input PHYEMAC0RXCHARISCOMMA;
    input PHYEMAC0RXCHARISK;
    input PHYEMAC0RXCHECKINGCRC;
    input PHYEMAC0RXCLK;
    input PHYEMAC0RXCOMMADET;
    input PHYEMAC0RXDISPERR;
    input PHYEMAC0RXDV;
    input PHYEMAC0RXER;
    input PHYEMAC0RXNOTINTABLE;
    input PHYEMAC0RXRUNDISP;
    input PHYEMAC0SIGNALDET;
    input PHYEMAC0TXBUFERR;
    input PHYEMAC0TXGMIIMIICLKIN;
    input PHYEMAC1COL;
    input PHYEMAC1CRS;
    input PHYEMAC1GTXCLK;
    input PHYEMAC1MCLKIN;
    input PHYEMAC1MDIN;
    input PHYEMAC1MIITXCLK;
    input PHYEMAC1RXBUFERR;
    input PHYEMAC1RXCHARISCOMMA;
    input PHYEMAC1RXCHARISK;
    input PHYEMAC1RXCHECKINGCRC;
    input PHYEMAC1RXCLK;
    input PHYEMAC1RXCOMMADET;
    input PHYEMAC1RXDISPERR;
    input PHYEMAC1RXDV;
    input PHYEMAC1RXER;
    input PHYEMAC1RXNOTINTABLE;
    input PHYEMAC1RXRUNDISP;
    input PHYEMAC1SIGNALDET;
    input PHYEMAC1TXBUFERR;
    input PHYEMAC1TXGMIIMIICLKIN;
    input RESET;
    input [0:31] DCREMACDBUS;
    input [0:9] DCREMACABUS;
    input [15:0] CLIENTEMAC0PAUSEVAL;
    input [15:0] CLIENTEMAC0TXD;
    input [15:0] CLIENTEMAC1PAUSEVAL;
    input [15:0] CLIENTEMAC1TXD;
    input [1:0] HOSTOPCODE;
    input [1:0] PHYEMAC0RXBUFSTATUS;
    input [1:0] PHYEMAC0RXLOSSOFSYNC;
    input [1:0] PHYEMAC1RXBUFSTATUS;
    input [1:0] PHYEMAC1RXLOSSOFSYNC;
    input [2:0] PHYEMAC0RXCLKCORCNT;
    input [2:0] PHYEMAC1RXCLKCORCNT;
    input [31:0] HOSTWRDATA;
    input [4:0] PHYEMAC0PHYAD;
    input [4:0] PHYEMAC1PHYAD;
    input [7:0] CLIENTEMAC0TXIFGDELAY;
    input [7:0] CLIENTEMAC1TXIFGDELAY;
    input [7:0] PHYEMAC0RXD;
    input [7:0] PHYEMAC1RXD;
    input [9:0] HOSTADDR;
endmodule

module TEMAC_SINGLE (...);
    parameter EMAC_1000BASEX_ENABLE = "FALSE";
    parameter EMAC_ADDRFILTER_ENABLE = "FALSE";
    parameter EMAC_BYTEPHY = "FALSE";
    parameter EMAC_CTRLLENCHECK_DISABLE = "FALSE";
    parameter [0:7] EMAC_DCRBASEADDR = 8'h00;
    parameter EMAC_GTLOOPBACK = "FALSE";
    parameter EMAC_HOST_ENABLE = "FALSE";
    parameter [8:0] EMAC_LINKTIMERVAL = 9'h000;
    parameter EMAC_LTCHECK_DISABLE = "FALSE";
    parameter EMAC_MDIO_ENABLE = "FALSE";
    parameter EMAC_MDIO_IGNORE_PHYADZERO = "FALSE";
    parameter [47:0] EMAC_PAUSEADDR = 48'h000000000000;
    parameter EMAC_PHYINITAUTONEG_ENABLE = "FALSE";
    parameter EMAC_PHYISOLATE = "FALSE";
    parameter EMAC_PHYLOOPBACKMSB = "FALSE";
    parameter EMAC_PHYPOWERDOWN = "FALSE";
    parameter EMAC_PHYRESET = "FALSE";
    parameter EMAC_RGMII_ENABLE = "FALSE";
    parameter EMAC_RX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC_RXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC_RXHALFDUPLEX = "FALSE";
    parameter EMAC_RXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC_RXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC_RXRESET = "FALSE";
    parameter EMAC_RXVLAN_ENABLE = "FALSE";
    parameter EMAC_RX_ENABLE = "TRUE";
    parameter EMAC_SGMII_ENABLE = "FALSE";
    parameter EMAC_SPEED_LSB = "FALSE";
    parameter EMAC_SPEED_MSB = "FALSE";
    parameter EMAC_TX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC_TXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC_TXHALFDUPLEX = "FALSE";
    parameter EMAC_TXIFGADJUST_ENABLE = "FALSE";
    parameter EMAC_TXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC_TXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC_TXRESET = "FALSE";
    parameter EMAC_TXVLAN_ENABLE = "FALSE";
    parameter EMAC_TX_ENABLE = "TRUE";
    parameter [47:0] EMAC_UNICASTADDR = 48'h000000000000;
    parameter EMAC_UNIDIRECTION_ENABLE = "FALSE";
    parameter EMAC_USECLKEN = "FALSE";
    parameter SIM_VERSION = "1.0";
    output DCRHOSTDONEIR;
    output EMACCLIENTANINTERRUPT;
    output EMACCLIENTRXBADFRAME;
    output EMACCLIENTRXCLIENTCLKOUT;
    output EMACCLIENTRXDVLD;
    output EMACCLIENTRXDVLDMSW;
    output EMACCLIENTRXFRAMEDROP;
    output EMACCLIENTRXGOODFRAME;
    output EMACCLIENTRXSTATSBYTEVLD;
    output EMACCLIENTRXSTATSVLD;
    output EMACCLIENTTXACK;
    output EMACCLIENTTXCLIENTCLKOUT;
    output EMACCLIENTTXCOLLISION;
    output EMACCLIENTTXRETRANSMIT;
    output EMACCLIENTTXSTATS;
    output EMACCLIENTTXSTATSBYTEVLD;
    output EMACCLIENTTXSTATSVLD;
    output EMACDCRACK;
    output EMACPHYENCOMMAALIGN;
    output EMACPHYLOOPBACKMSB;
    output EMACPHYMCLKOUT;
    output EMACPHYMDOUT;
    output EMACPHYMDTRI;
    output EMACPHYMGTRXRESET;
    output EMACPHYMGTTXRESET;
    output EMACPHYPOWERDOWN;
    output EMACPHYSYNCACQSTATUS;
    output EMACPHYTXCHARDISPMODE;
    output EMACPHYTXCHARDISPVAL;
    output EMACPHYTXCHARISK;
    output EMACPHYTXCLK;
    output EMACPHYTXEN;
    output EMACPHYTXER;
    output EMACPHYTXGMIIMIICLKOUT;
    output EMACSPEEDIS10100;
    output HOSTMIIMRDY;
    output [0:31] EMACDCRDBUS;
    output [15:0] EMACCLIENTRXD;
    output [31:0] HOSTRDDATA;
    output [6:0] EMACCLIENTRXSTATS;
    output [7:0] EMACPHYTXD;
    input CLIENTEMACDCMLOCKED;
    input CLIENTEMACPAUSEREQ;
    input CLIENTEMACRXCLIENTCLKIN;
    input CLIENTEMACTXCLIENTCLKIN;
    input CLIENTEMACTXDVLD;
    input CLIENTEMACTXDVLDMSW;
    input CLIENTEMACTXFIRSTBYTE;
    input CLIENTEMACTXUNDERRUN;
    input DCREMACCLK;
    input DCREMACENABLE;
    input DCREMACREAD;
    input DCREMACWRITE;
    input HOSTCLK;
    input HOSTMIIMSEL;
    input HOSTREQ;
    input PHYEMACCOL;
    input PHYEMACCRS;
    input PHYEMACGTXCLK;
    input PHYEMACMCLKIN;
    input PHYEMACMDIN;
    input PHYEMACMIITXCLK;
    input PHYEMACRXCHARISCOMMA;
    input PHYEMACRXCHARISK;
    input PHYEMACRXCLK;
    input PHYEMACRXDISPERR;
    input PHYEMACRXDV;
    input PHYEMACRXER;
    input PHYEMACRXNOTINTABLE;
    input PHYEMACRXRUNDISP;
    input PHYEMACSIGNALDET;
    input PHYEMACTXBUFERR;
    input PHYEMACTXGMIIMIICLKIN;
    input RESET;
    input [0:31] DCREMACDBUS;
    input [0:9] DCREMACABUS;
    input [15:0] CLIENTEMACPAUSEVAL;
    input [15:0] CLIENTEMACTXD;
    input [1:0] HOSTOPCODE;
    input [1:0] PHYEMACRXBUFSTATUS;
    input [2:0] PHYEMACRXCLKCORCNT;
    input [31:0] HOSTWRDATA;
    input [4:0] PHYEMACPHYAD;
    input [7:0] CLIENTEMACTXIFGDELAY;
    input [7:0] PHYEMACRXD;
    input [9:0] HOSTADDR;
endmodule

module CMAC (...);
    parameter CTL_PTP_TRANSPCLK_MODE = "FALSE";
    parameter CTL_RX_CHECK_ACK = "TRUE";
    parameter CTL_RX_CHECK_PREAMBLE = "FALSE";
    parameter CTL_RX_CHECK_SFD = "FALSE";
    parameter CTL_RX_DELETE_FCS = "TRUE";
    parameter [15:0] CTL_RX_ETYPE_GCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_GPP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PPP = 16'h8808;
    parameter CTL_RX_FORWARD_CONTROL = "FALSE";
    parameter CTL_RX_IGNORE_FCS = "FALSE";
    parameter [14:0] CTL_RX_MAX_PACKET_LEN = 15'h2580;
    parameter [7:0] CTL_RX_MIN_PACKET_LEN = 8'h40;
    parameter [15:0] CTL_RX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_RX_OPCODE_MAX_GCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MAX_PCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MIN_GCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_MIN_PCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_PPP = 16'h0001;
    parameter [47:0] CTL_RX_PAUSE_DA_MCAST = 48'h0180C2000001;
    parameter [47:0] CTL_RX_PAUSE_DA_UCAST = 48'h000000000000;
    parameter [47:0] CTL_RX_PAUSE_SA = 48'h000000000000;
    parameter CTL_RX_PROCESS_LFI = "FALSE";
    parameter [15:0] CTL_RX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_RX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_RX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_RX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_RX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_RX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_RX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_RX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_RX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_RX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_RX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_RX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_RX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_RX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_RX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_RX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_RX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_RX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_RX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [47:0] CTL_TX_DA_GPP = 48'h0180C2000001;
    parameter [47:0] CTL_TX_DA_PPP = 48'h0180C2000001;
    parameter [15:0] CTL_TX_ETHERTYPE_GPP = 16'h8808;
    parameter [15:0] CTL_TX_ETHERTYPE_PPP = 16'h8808;
    parameter CTL_TX_FCS_INS_ENABLE = "TRUE";
    parameter CTL_TX_IGNORE_FCS = "FALSE";
    parameter [15:0] CTL_TX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_TX_OPCODE_PPP = 16'h0001;
    parameter CTL_TX_PTP_1STEP_ENABLE = "FALSE";
    parameter [10:0] CTL_TX_PTP_LATENCY_ADJUST = 11'h2C1;
    parameter [47:0] CTL_TX_SA_GPP = 48'h000000000000;
    parameter [47:0] CTL_TX_SA_PPP = 48'h000000000000;
    parameter [15:0] CTL_TX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_TX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_TX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_TX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_TX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_TX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_TX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_TX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_TX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_TX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_TX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_TX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_TX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_TX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_TX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_TX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_TX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_TX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_TX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter SIM_VERSION = "2.0";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [6:0] RX_LANE_ALIGNER_FILL_0;
    output [6:0] RX_LANE_ALIGNER_FILL_1;
    output [6:0] RX_LANE_ALIGNER_FILL_10;
    output [6:0] RX_LANE_ALIGNER_FILL_11;
    output [6:0] RX_LANE_ALIGNER_FILL_12;
    output [6:0] RX_LANE_ALIGNER_FILL_13;
    output [6:0] RX_LANE_ALIGNER_FILL_14;
    output [6:0] RX_LANE_ALIGNER_FILL_15;
    output [6:0] RX_LANE_ALIGNER_FILL_16;
    output [6:0] RX_LANE_ALIGNER_FILL_17;
    output [6:0] RX_LANE_ALIGNER_FILL_18;
    output [6:0] RX_LANE_ALIGNER_FILL_19;
    output [6:0] RX_LANE_ALIGNER_FILL_2;
    output [6:0] RX_LANE_ALIGNER_FILL_3;
    output [6:0] RX_LANE_ALIGNER_FILL_4;
    output [6:0] RX_LANE_ALIGNER_FILL_5;
    output [6:0] RX_LANE_ALIGNER_FILL_6;
    output [6:0] RX_LANE_ALIGNER_FILL_7;
    output [6:0] RX_LANE_ALIGNER_FILL_8;
    output [6:0] RX_LANE_ALIGNER_FILL_9;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output [4:0] RX_PTP_PCSLANE_OUT;
    output [79:0] RX_PTP_TSTAMP_OUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [6:0] STAT_RX_BAD_CODE;
    output [3:0] STAT_RX_BAD_FCS;
    output STAT_RX_BAD_PREAMBLE;
    output STAT_RX_BAD_SFD;
    output STAT_RX_BIP_ERR_0;
    output STAT_RX_BIP_ERR_1;
    output STAT_RX_BIP_ERR_10;
    output STAT_RX_BIP_ERR_11;
    output STAT_RX_BIP_ERR_12;
    output STAT_RX_BIP_ERR_13;
    output STAT_RX_BIP_ERR_14;
    output STAT_RX_BIP_ERR_15;
    output STAT_RX_BIP_ERR_16;
    output STAT_RX_BIP_ERR_17;
    output STAT_RX_BIP_ERR_18;
    output STAT_RX_BIP_ERR_19;
    output STAT_RX_BIP_ERR_2;
    output STAT_RX_BIP_ERR_3;
    output STAT_RX_BIP_ERR_4;
    output STAT_RX_BIP_ERR_5;
    output STAT_RX_BIP_ERR_6;
    output STAT_RX_BIP_ERR_7;
    output STAT_RX_BIP_ERR_8;
    output STAT_RX_BIP_ERR_9;
    output [19:0] STAT_RX_BLOCK_LOCK;
    output STAT_RX_BROADCAST;
    output [3:0] STAT_RX_FRAGMENT;
    output [3:0] STAT_RX_FRAMING_ERR_0;
    output [3:0] STAT_RX_FRAMING_ERR_1;
    output [3:0] STAT_RX_FRAMING_ERR_10;
    output [3:0] STAT_RX_FRAMING_ERR_11;
    output [3:0] STAT_RX_FRAMING_ERR_12;
    output [3:0] STAT_RX_FRAMING_ERR_13;
    output [3:0] STAT_RX_FRAMING_ERR_14;
    output [3:0] STAT_RX_FRAMING_ERR_15;
    output [3:0] STAT_RX_FRAMING_ERR_16;
    output [3:0] STAT_RX_FRAMING_ERR_17;
    output [3:0] STAT_RX_FRAMING_ERR_18;
    output [3:0] STAT_RX_FRAMING_ERR_19;
    output [3:0] STAT_RX_FRAMING_ERR_2;
    output [3:0] STAT_RX_FRAMING_ERR_3;
    output [3:0] STAT_RX_FRAMING_ERR_4;
    output [3:0] STAT_RX_FRAMING_ERR_5;
    output [3:0] STAT_RX_FRAMING_ERR_6;
    output [3:0] STAT_RX_FRAMING_ERR_7;
    output [3:0] STAT_RX_FRAMING_ERR_8;
    output [3:0] STAT_RX_FRAMING_ERR_9;
    output STAT_RX_FRAMING_ERR_VALID_0;
    output STAT_RX_FRAMING_ERR_VALID_1;
    output STAT_RX_FRAMING_ERR_VALID_10;
    output STAT_RX_FRAMING_ERR_VALID_11;
    output STAT_RX_FRAMING_ERR_VALID_12;
    output STAT_RX_FRAMING_ERR_VALID_13;
    output STAT_RX_FRAMING_ERR_VALID_14;
    output STAT_RX_FRAMING_ERR_VALID_15;
    output STAT_RX_FRAMING_ERR_VALID_16;
    output STAT_RX_FRAMING_ERR_VALID_17;
    output STAT_RX_FRAMING_ERR_VALID_18;
    output STAT_RX_FRAMING_ERR_VALID_19;
    output STAT_RX_FRAMING_ERR_VALID_2;
    output STAT_RX_FRAMING_ERR_VALID_3;
    output STAT_RX_FRAMING_ERR_VALID_4;
    output STAT_RX_FRAMING_ERR_VALID_5;
    output STAT_RX_FRAMING_ERR_VALID_6;
    output STAT_RX_FRAMING_ERR_VALID_7;
    output STAT_RX_FRAMING_ERR_VALID_8;
    output STAT_RX_FRAMING_ERR_VALID_9;
    output STAT_RX_GOT_SIGNAL_OS;
    output STAT_RX_HI_BER;
    output STAT_RX_INRANGEERR;
    output STAT_RX_INTERNAL_LOCAL_FAULT;
    output STAT_RX_JABBER;
    output [7:0] STAT_RX_LANE0_VLM_BIP7;
    output STAT_RX_LANE0_VLM_BIP7_VALID;
    output STAT_RX_LOCAL_FAULT;
    output [19:0] STAT_RX_MF_ERR;
    output [19:0] STAT_RX_MF_LEN_ERR;
    output [19:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MULTICAST;
    output STAT_RX_OVERSIZE;
    output STAT_RX_PACKET_1024_1518_BYTES;
    output STAT_RX_PACKET_128_255_BYTES;
    output STAT_RX_PACKET_1519_1522_BYTES;
    output STAT_RX_PACKET_1523_1548_BYTES;
    output STAT_RX_PACKET_1549_2047_BYTES;
    output STAT_RX_PACKET_2048_4095_BYTES;
    output STAT_RX_PACKET_256_511_BYTES;
    output STAT_RX_PACKET_4096_8191_BYTES;
    output STAT_RX_PACKET_512_1023_BYTES;
    output STAT_RX_PACKET_64_BYTES;
    output STAT_RX_PACKET_65_127_BYTES;
    output STAT_RX_PACKET_8192_9215_BYTES;
    output STAT_RX_PACKET_BAD_FCS;
    output STAT_RX_PACKET_LARGE;
    output [3:0] STAT_RX_PACKET_SMALL;
    output STAT_RX_PAUSE;
    output [15:0] STAT_RX_PAUSE_QUANTA0;
    output [15:0] STAT_RX_PAUSE_QUANTA1;
    output [15:0] STAT_RX_PAUSE_QUANTA2;
    output [15:0] STAT_RX_PAUSE_QUANTA3;
    output [15:0] STAT_RX_PAUSE_QUANTA4;
    output [15:0] STAT_RX_PAUSE_QUANTA5;
    output [15:0] STAT_RX_PAUSE_QUANTA6;
    output [15:0] STAT_RX_PAUSE_QUANTA7;
    output [15:0] STAT_RX_PAUSE_QUANTA8;
    output [8:0] STAT_RX_PAUSE_REQ;
    output [8:0] STAT_RX_PAUSE_VALID;
    output STAT_RX_RECEIVED_LOCAL_FAULT;
    output STAT_RX_REMOTE_FAULT;
    output STAT_RX_STATUS;
    output [3:0] STAT_RX_STOMPED_FCS;
    output [19:0] STAT_RX_SYNCED;
    output [19:0] STAT_RX_SYNCED_ERR;
    output [2:0] STAT_RX_TEST_PATTERN_MISMATCH;
    output STAT_RX_TOOLONG;
    output [7:0] STAT_RX_TOTAL_BYTES;
    output [13:0] STAT_RX_TOTAL_GOOD_BYTES;
    output STAT_RX_TOTAL_GOOD_PACKETS;
    output [3:0] STAT_RX_TOTAL_PACKETS;
    output STAT_RX_TRUNCATED;
    output [3:0] STAT_RX_UNDERSIZE;
    output STAT_RX_UNICAST;
    output STAT_RX_USER_PAUSE;
    output STAT_RX_VLAN;
    output [19:0] STAT_RX_VL_DEMUXED;
    output [4:0] STAT_RX_VL_NUMBER_0;
    output [4:0] STAT_RX_VL_NUMBER_1;
    output [4:0] STAT_RX_VL_NUMBER_10;
    output [4:0] STAT_RX_VL_NUMBER_11;
    output [4:0] STAT_RX_VL_NUMBER_12;
    output [4:0] STAT_RX_VL_NUMBER_13;
    output [4:0] STAT_RX_VL_NUMBER_14;
    output [4:0] STAT_RX_VL_NUMBER_15;
    output [4:0] STAT_RX_VL_NUMBER_16;
    output [4:0] STAT_RX_VL_NUMBER_17;
    output [4:0] STAT_RX_VL_NUMBER_18;
    output [4:0] STAT_RX_VL_NUMBER_19;
    output [4:0] STAT_RX_VL_NUMBER_2;
    output [4:0] STAT_RX_VL_NUMBER_3;
    output [4:0] STAT_RX_VL_NUMBER_4;
    output [4:0] STAT_RX_VL_NUMBER_5;
    output [4:0] STAT_RX_VL_NUMBER_6;
    output [4:0] STAT_RX_VL_NUMBER_7;
    output [4:0] STAT_RX_VL_NUMBER_8;
    output [4:0] STAT_RX_VL_NUMBER_9;
    output STAT_TX_BAD_FCS;
    output STAT_TX_BROADCAST;
    output STAT_TX_FRAME_ERROR;
    output STAT_TX_LOCAL_FAULT;
    output STAT_TX_MULTICAST;
    output STAT_TX_PACKET_1024_1518_BYTES;
    output STAT_TX_PACKET_128_255_BYTES;
    output STAT_TX_PACKET_1519_1522_BYTES;
    output STAT_TX_PACKET_1523_1548_BYTES;
    output STAT_TX_PACKET_1549_2047_BYTES;
    output STAT_TX_PACKET_2048_4095_BYTES;
    output STAT_TX_PACKET_256_511_BYTES;
    output STAT_TX_PACKET_4096_8191_BYTES;
    output STAT_TX_PACKET_512_1023_BYTES;
    output STAT_TX_PACKET_64_BYTES;
    output STAT_TX_PACKET_65_127_BYTES;
    output STAT_TX_PACKET_8192_9215_BYTES;
    output STAT_TX_PACKET_LARGE;
    output STAT_TX_PACKET_SMALL;
    output STAT_TX_PAUSE;
    output [8:0] STAT_TX_PAUSE_VALID;
    output STAT_TX_PTP_FIFO_READ_ERROR;
    output STAT_TX_PTP_FIFO_WRITE_ERROR;
    output [6:0] STAT_TX_TOTAL_BYTES;
    output [13:0] STAT_TX_TOTAL_GOOD_BYTES;
    output STAT_TX_TOTAL_GOOD_PACKETS;
    output STAT_TX_TOTAL_PACKETS;
    output STAT_TX_UNICAST;
    output STAT_TX_USER_PAUSE;
    output STAT_TX_VLAN;
    output TX_OVFOUT;
    output [4:0] TX_PTP_PCSLANE_OUT;
    output [79:0] TX_PTP_TSTAMP_OUT;
    output [15:0] TX_PTP_TSTAMP_TAG_OUT;
    output TX_PTP_TSTAMP_VALID_OUT;
    output TX_RDYOUT;
    output [15:0] TX_SERDES_ALT_DATA0;
    output [15:0] TX_SERDES_ALT_DATA1;
    output [15:0] TX_SERDES_ALT_DATA2;
    output [15:0] TX_SERDES_ALT_DATA3;
    output [63:0] TX_SERDES_DATA0;
    output [63:0] TX_SERDES_DATA1;
    output [63:0] TX_SERDES_DATA2;
    output [63:0] TX_SERDES_DATA3;
    output [31:0] TX_SERDES_DATA4;
    output [31:0] TX_SERDES_DATA5;
    output [31:0] TX_SERDES_DATA6;
    output [31:0] TX_SERDES_DATA7;
    output [31:0] TX_SERDES_DATA8;
    output [31:0] TX_SERDES_DATA9;
    output TX_UNFOUT;
    input CTL_CAUI4_MODE;
    input CTL_RX_CHECK_ETYPE_GCP;
    input CTL_RX_CHECK_ETYPE_GPP;
    input CTL_RX_CHECK_ETYPE_PCP;
    input CTL_RX_CHECK_ETYPE_PPP;
    input CTL_RX_CHECK_MCAST_GCP;
    input CTL_RX_CHECK_MCAST_GPP;
    input CTL_RX_CHECK_MCAST_PCP;
    input CTL_RX_CHECK_MCAST_PPP;
    input CTL_RX_CHECK_OPCODE_GCP;
    input CTL_RX_CHECK_OPCODE_GPP;
    input CTL_RX_CHECK_OPCODE_PCP;
    input CTL_RX_CHECK_OPCODE_PPP;
    input CTL_RX_CHECK_SA_GCP;
    input CTL_RX_CHECK_SA_GPP;
    input CTL_RX_CHECK_SA_PCP;
    input CTL_RX_CHECK_SA_PPP;
    input CTL_RX_CHECK_UCAST_GCP;
    input CTL_RX_CHECK_UCAST_GPP;
    input CTL_RX_CHECK_UCAST_PCP;
    input CTL_RX_CHECK_UCAST_PPP;
    input CTL_RX_ENABLE;
    input CTL_RX_ENABLE_GCP;
    input CTL_RX_ENABLE_GPP;
    input CTL_RX_ENABLE_PCP;
    input CTL_RX_ENABLE_PPP;
    input CTL_RX_FORCE_RESYNC;
    input [8:0] CTL_RX_PAUSE_ACK;
    input [8:0] CTL_RX_PAUSE_ENABLE;
    input [79:0] CTL_RX_SYSTEMTIMERIN;
    input CTL_RX_TEST_PATTERN;
    input CTL_TX_ENABLE;
    input CTL_TX_LANE0_VLM_BIP7_OVERRIDE;
    input [7:0] CTL_TX_LANE0_VLM_BIP7_OVERRIDE_VALUE;
    input [8:0] CTL_TX_PAUSE_ENABLE;
    input [15:0] CTL_TX_PAUSE_QUANTA0;
    input [15:0] CTL_TX_PAUSE_QUANTA1;
    input [15:0] CTL_TX_PAUSE_QUANTA2;
    input [15:0] CTL_TX_PAUSE_QUANTA3;
    input [15:0] CTL_TX_PAUSE_QUANTA4;
    input [15:0] CTL_TX_PAUSE_QUANTA5;
    input [15:0] CTL_TX_PAUSE_QUANTA6;
    input [15:0] CTL_TX_PAUSE_QUANTA7;
    input [15:0] CTL_TX_PAUSE_QUANTA8;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER0;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER1;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER2;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER3;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER4;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER5;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER6;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER7;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER8;
    input [8:0] CTL_TX_PAUSE_REQ;
    input CTL_TX_PTP_VLANE_ADJUST_MODE;
    input CTL_TX_RESEND_PAUSE;
    input CTL_TX_SEND_IDLE;
    input CTL_TX_SEND_RFI;
    input [79:0] CTL_TX_SYSTEMTIMERIN;
    input CTL_TX_TEST_PATTERN;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input RX_CLK;
    input RX_RESET;
    input [15:0] RX_SERDES_ALT_DATA0;
    input [15:0] RX_SERDES_ALT_DATA1;
    input [15:0] RX_SERDES_ALT_DATA2;
    input [15:0] RX_SERDES_ALT_DATA3;
    input [9:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA0;
    input [63:0] RX_SERDES_DATA1;
    input [63:0] RX_SERDES_DATA2;
    input [63:0] RX_SERDES_DATA3;
    input [31:0] RX_SERDES_DATA4;
    input [31:0] RX_SERDES_DATA5;
    input [31:0] RX_SERDES_DATA6;
    input [31:0] RX_SERDES_DATA7;
    input [31:0] RX_SERDES_DATA8;
    input [31:0] RX_SERDES_DATA9;
    input [9:0] RX_SERDES_RESET;
    input TX_CLK;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input [1:0] TX_PTP_1588OP_IN;
    input [15:0] TX_PTP_CHKSUM_OFFSET_IN;
    input [63:0] TX_PTP_RXTSTAMP_IN;
    input [15:0] TX_PTP_TAG_FIELD_IN;
    input [15:0] TX_PTP_TSTAMP_OFFSET_IN;
    input TX_PTP_UPD_CHKSUM_IN;
    input TX_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module CMACE4 (...);
    parameter CTL_PTP_TRANSPCLK_MODE = "FALSE";
    parameter CTL_RX_CHECK_ACK = "TRUE";
    parameter CTL_RX_CHECK_PREAMBLE = "FALSE";
    parameter CTL_RX_CHECK_SFD = "FALSE";
    parameter CTL_RX_DELETE_FCS = "TRUE";
    parameter [15:0] CTL_RX_ETYPE_GCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_GPP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PPP = 16'h8808;
    parameter CTL_RX_FORWARD_CONTROL = "FALSE";
    parameter CTL_RX_IGNORE_FCS = "FALSE";
    parameter [14:0] CTL_RX_MAX_PACKET_LEN = 15'h2580;
    parameter [7:0] CTL_RX_MIN_PACKET_LEN = 8'h40;
    parameter [15:0] CTL_RX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_RX_OPCODE_MAX_GCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MAX_PCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MIN_GCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_MIN_PCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_PPP = 16'h0001;
    parameter [47:0] CTL_RX_PAUSE_DA_MCAST = 48'h0180C2000001;
    parameter [47:0] CTL_RX_PAUSE_DA_UCAST = 48'h000000000000;
    parameter [47:0] CTL_RX_PAUSE_SA = 48'h000000000000;
    parameter CTL_RX_PROCESS_LFI = "FALSE";
    parameter [8:0] CTL_RX_RSFEC_AM_THRESHOLD = 9'h046;
    parameter [1:0] CTL_RX_RSFEC_FILL_ADJUST = 2'h0;
    parameter [15:0] CTL_RX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_RX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_RX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_RX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_RX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_RX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_RX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_RX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_RX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_RX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_RX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_RX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_RX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_RX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_RX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_RX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_RX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_RX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_RX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter CTL_TX_CUSTOM_PREAMBLE_ENABLE = "FALSE";
    parameter [47:0] CTL_TX_DA_GPP = 48'h0180C2000001;
    parameter [47:0] CTL_TX_DA_PPP = 48'h0180C2000001;
    parameter [15:0] CTL_TX_ETHERTYPE_GPP = 16'h8808;
    parameter [15:0] CTL_TX_ETHERTYPE_PPP = 16'h8808;
    parameter CTL_TX_FCS_INS_ENABLE = "TRUE";
    parameter CTL_TX_IGNORE_FCS = "FALSE";
    parameter [3:0] CTL_TX_IPG_VALUE = 4'hC;
    parameter [15:0] CTL_TX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_TX_OPCODE_PPP = 16'h0001;
    parameter CTL_TX_PTP_1STEP_ENABLE = "FALSE";
    parameter [10:0] CTL_TX_PTP_LATENCY_ADJUST = 11'h2C1;
    parameter [47:0] CTL_TX_SA_GPP = 48'h000000000000;
    parameter [47:0] CTL_TX_SA_PPP = 48'h000000000000;
    parameter [15:0] CTL_TX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_TX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_TX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_TX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_TX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_TX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_TX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_TX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_TX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_TX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_TX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_TX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_TX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_TX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_TX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_TX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_TX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_TX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_TX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [329:0] RSFEC_BYPASS_RX_DOUT;
    output RSFEC_BYPASS_RX_DOUT_CW_START;
    output RSFEC_BYPASS_RX_DOUT_VALID;
    output [329:0] RSFEC_BYPASS_TX_DOUT;
    output RSFEC_BYPASS_TX_DOUT_CW_START;
    output RSFEC_BYPASS_TX_DOUT_VALID;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [6:0] RX_LANE_ALIGNER_FILL_0;
    output [6:0] RX_LANE_ALIGNER_FILL_1;
    output [6:0] RX_LANE_ALIGNER_FILL_10;
    output [6:0] RX_LANE_ALIGNER_FILL_11;
    output [6:0] RX_LANE_ALIGNER_FILL_12;
    output [6:0] RX_LANE_ALIGNER_FILL_13;
    output [6:0] RX_LANE_ALIGNER_FILL_14;
    output [6:0] RX_LANE_ALIGNER_FILL_15;
    output [6:0] RX_LANE_ALIGNER_FILL_16;
    output [6:0] RX_LANE_ALIGNER_FILL_17;
    output [6:0] RX_LANE_ALIGNER_FILL_18;
    output [6:0] RX_LANE_ALIGNER_FILL_19;
    output [6:0] RX_LANE_ALIGNER_FILL_2;
    output [6:0] RX_LANE_ALIGNER_FILL_3;
    output [6:0] RX_LANE_ALIGNER_FILL_4;
    output [6:0] RX_LANE_ALIGNER_FILL_5;
    output [6:0] RX_LANE_ALIGNER_FILL_6;
    output [6:0] RX_LANE_ALIGNER_FILL_7;
    output [6:0] RX_LANE_ALIGNER_FILL_8;
    output [6:0] RX_LANE_ALIGNER_FILL_9;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output [7:0] RX_OTN_BIP8_0;
    output [7:0] RX_OTN_BIP8_1;
    output [7:0] RX_OTN_BIP8_2;
    output [7:0] RX_OTN_BIP8_3;
    output [7:0] RX_OTN_BIP8_4;
    output [65:0] RX_OTN_DATA_0;
    output [65:0] RX_OTN_DATA_1;
    output [65:0] RX_OTN_DATA_2;
    output [65:0] RX_OTN_DATA_3;
    output [65:0] RX_OTN_DATA_4;
    output RX_OTN_ENA;
    output RX_OTN_LANE0;
    output RX_OTN_VLMARKER;
    output [55:0] RX_PREOUT;
    output [4:0] RX_PTP_PCSLANE_OUT;
    output [79:0] RX_PTP_TSTAMP_OUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [2:0] STAT_RX_BAD_CODE;
    output [2:0] STAT_RX_BAD_FCS;
    output STAT_RX_BAD_PREAMBLE;
    output STAT_RX_BAD_SFD;
    output STAT_RX_BIP_ERR_0;
    output STAT_RX_BIP_ERR_1;
    output STAT_RX_BIP_ERR_10;
    output STAT_RX_BIP_ERR_11;
    output STAT_RX_BIP_ERR_12;
    output STAT_RX_BIP_ERR_13;
    output STAT_RX_BIP_ERR_14;
    output STAT_RX_BIP_ERR_15;
    output STAT_RX_BIP_ERR_16;
    output STAT_RX_BIP_ERR_17;
    output STAT_RX_BIP_ERR_18;
    output STAT_RX_BIP_ERR_19;
    output STAT_RX_BIP_ERR_2;
    output STAT_RX_BIP_ERR_3;
    output STAT_RX_BIP_ERR_4;
    output STAT_RX_BIP_ERR_5;
    output STAT_RX_BIP_ERR_6;
    output STAT_RX_BIP_ERR_7;
    output STAT_RX_BIP_ERR_8;
    output STAT_RX_BIP_ERR_9;
    output [19:0] STAT_RX_BLOCK_LOCK;
    output STAT_RX_BROADCAST;
    output [2:0] STAT_RX_FRAGMENT;
    output [1:0] STAT_RX_FRAMING_ERR_0;
    output [1:0] STAT_RX_FRAMING_ERR_1;
    output [1:0] STAT_RX_FRAMING_ERR_10;
    output [1:0] STAT_RX_FRAMING_ERR_11;
    output [1:0] STAT_RX_FRAMING_ERR_12;
    output [1:0] STAT_RX_FRAMING_ERR_13;
    output [1:0] STAT_RX_FRAMING_ERR_14;
    output [1:0] STAT_RX_FRAMING_ERR_15;
    output [1:0] STAT_RX_FRAMING_ERR_16;
    output [1:0] STAT_RX_FRAMING_ERR_17;
    output [1:0] STAT_RX_FRAMING_ERR_18;
    output [1:0] STAT_RX_FRAMING_ERR_19;
    output [1:0] STAT_RX_FRAMING_ERR_2;
    output [1:0] STAT_RX_FRAMING_ERR_3;
    output [1:0] STAT_RX_FRAMING_ERR_4;
    output [1:0] STAT_RX_FRAMING_ERR_5;
    output [1:0] STAT_RX_FRAMING_ERR_6;
    output [1:0] STAT_RX_FRAMING_ERR_7;
    output [1:0] STAT_RX_FRAMING_ERR_8;
    output [1:0] STAT_RX_FRAMING_ERR_9;
    output STAT_RX_FRAMING_ERR_VALID_0;
    output STAT_RX_FRAMING_ERR_VALID_1;
    output STAT_RX_FRAMING_ERR_VALID_10;
    output STAT_RX_FRAMING_ERR_VALID_11;
    output STAT_RX_FRAMING_ERR_VALID_12;
    output STAT_RX_FRAMING_ERR_VALID_13;
    output STAT_RX_FRAMING_ERR_VALID_14;
    output STAT_RX_FRAMING_ERR_VALID_15;
    output STAT_RX_FRAMING_ERR_VALID_16;
    output STAT_RX_FRAMING_ERR_VALID_17;
    output STAT_RX_FRAMING_ERR_VALID_18;
    output STAT_RX_FRAMING_ERR_VALID_19;
    output STAT_RX_FRAMING_ERR_VALID_2;
    output STAT_RX_FRAMING_ERR_VALID_3;
    output STAT_RX_FRAMING_ERR_VALID_4;
    output STAT_RX_FRAMING_ERR_VALID_5;
    output STAT_RX_FRAMING_ERR_VALID_6;
    output STAT_RX_FRAMING_ERR_VALID_7;
    output STAT_RX_FRAMING_ERR_VALID_8;
    output STAT_RX_FRAMING_ERR_VALID_9;
    output STAT_RX_GOT_SIGNAL_OS;
    output STAT_RX_HI_BER;
    output STAT_RX_INRANGEERR;
    output STAT_RX_INTERNAL_LOCAL_FAULT;
    output STAT_RX_JABBER;
    output [7:0] STAT_RX_LANE0_VLM_BIP7;
    output STAT_RX_LANE0_VLM_BIP7_VALID;
    output STAT_RX_LOCAL_FAULT;
    output [19:0] STAT_RX_MF_ERR;
    output [19:0] STAT_RX_MF_LEN_ERR;
    output [19:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MULTICAST;
    output STAT_RX_OVERSIZE;
    output STAT_RX_PACKET_1024_1518_BYTES;
    output STAT_RX_PACKET_128_255_BYTES;
    output STAT_RX_PACKET_1519_1522_BYTES;
    output STAT_RX_PACKET_1523_1548_BYTES;
    output STAT_RX_PACKET_1549_2047_BYTES;
    output STAT_RX_PACKET_2048_4095_BYTES;
    output STAT_RX_PACKET_256_511_BYTES;
    output STAT_RX_PACKET_4096_8191_BYTES;
    output STAT_RX_PACKET_512_1023_BYTES;
    output STAT_RX_PACKET_64_BYTES;
    output STAT_RX_PACKET_65_127_BYTES;
    output STAT_RX_PACKET_8192_9215_BYTES;
    output STAT_RX_PACKET_BAD_FCS;
    output STAT_RX_PACKET_LARGE;
    output [2:0] STAT_RX_PACKET_SMALL;
    output STAT_RX_PAUSE;
    output [15:0] STAT_RX_PAUSE_QUANTA0;
    output [15:0] STAT_RX_PAUSE_QUANTA1;
    output [15:0] STAT_RX_PAUSE_QUANTA2;
    output [15:0] STAT_RX_PAUSE_QUANTA3;
    output [15:0] STAT_RX_PAUSE_QUANTA4;
    output [15:0] STAT_RX_PAUSE_QUANTA5;
    output [15:0] STAT_RX_PAUSE_QUANTA6;
    output [15:0] STAT_RX_PAUSE_QUANTA7;
    output [15:0] STAT_RX_PAUSE_QUANTA8;
    output [8:0] STAT_RX_PAUSE_REQ;
    output [8:0] STAT_RX_PAUSE_VALID;
    output STAT_RX_RECEIVED_LOCAL_FAULT;
    output STAT_RX_REMOTE_FAULT;
    output STAT_RX_RSFEC_AM_LOCK0;
    output STAT_RX_RSFEC_AM_LOCK1;
    output STAT_RX_RSFEC_AM_LOCK2;
    output STAT_RX_RSFEC_AM_LOCK3;
    output STAT_RX_RSFEC_CORRECTED_CW_INC;
    output STAT_RX_RSFEC_CW_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT0_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT1_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT2_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT3_INC;
    output STAT_RX_RSFEC_HI_SER;
    output STAT_RX_RSFEC_LANE_ALIGNMENT_STATUS;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_0;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_1;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_2;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_3;
    output [7:0] STAT_RX_RSFEC_LANE_MAPPING;
    output [31:0] STAT_RX_RSFEC_RSVD;
    output STAT_RX_RSFEC_UNCORRECTED_CW_INC;
    output STAT_RX_STATUS;
    output [2:0] STAT_RX_STOMPED_FCS;
    output [19:0] STAT_RX_SYNCED;
    output [19:0] STAT_RX_SYNCED_ERR;
    output [2:0] STAT_RX_TEST_PATTERN_MISMATCH;
    output STAT_RX_TOOLONG;
    output [6:0] STAT_RX_TOTAL_BYTES;
    output [13:0] STAT_RX_TOTAL_GOOD_BYTES;
    output STAT_RX_TOTAL_GOOD_PACKETS;
    output [2:0] STAT_RX_TOTAL_PACKETS;
    output STAT_RX_TRUNCATED;
    output [2:0] STAT_RX_UNDERSIZE;
    output STAT_RX_UNICAST;
    output STAT_RX_USER_PAUSE;
    output STAT_RX_VLAN;
    output [19:0] STAT_RX_VL_DEMUXED;
    output [4:0] STAT_RX_VL_NUMBER_0;
    output [4:0] STAT_RX_VL_NUMBER_1;
    output [4:0] STAT_RX_VL_NUMBER_10;
    output [4:0] STAT_RX_VL_NUMBER_11;
    output [4:0] STAT_RX_VL_NUMBER_12;
    output [4:0] STAT_RX_VL_NUMBER_13;
    output [4:0] STAT_RX_VL_NUMBER_14;
    output [4:0] STAT_RX_VL_NUMBER_15;
    output [4:0] STAT_RX_VL_NUMBER_16;
    output [4:0] STAT_RX_VL_NUMBER_17;
    output [4:0] STAT_RX_VL_NUMBER_18;
    output [4:0] STAT_RX_VL_NUMBER_19;
    output [4:0] STAT_RX_VL_NUMBER_2;
    output [4:0] STAT_RX_VL_NUMBER_3;
    output [4:0] STAT_RX_VL_NUMBER_4;
    output [4:0] STAT_RX_VL_NUMBER_5;
    output [4:0] STAT_RX_VL_NUMBER_6;
    output [4:0] STAT_RX_VL_NUMBER_7;
    output [4:0] STAT_RX_VL_NUMBER_8;
    output [4:0] STAT_RX_VL_NUMBER_9;
    output STAT_TX_BAD_FCS;
    output STAT_TX_BROADCAST;
    output STAT_TX_FRAME_ERROR;
    output STAT_TX_LOCAL_FAULT;
    output STAT_TX_MULTICAST;
    output STAT_TX_PACKET_1024_1518_BYTES;
    output STAT_TX_PACKET_128_255_BYTES;
    output STAT_TX_PACKET_1519_1522_BYTES;
    output STAT_TX_PACKET_1523_1548_BYTES;
    output STAT_TX_PACKET_1549_2047_BYTES;
    output STAT_TX_PACKET_2048_4095_BYTES;
    output STAT_TX_PACKET_256_511_BYTES;
    output STAT_TX_PACKET_4096_8191_BYTES;
    output STAT_TX_PACKET_512_1023_BYTES;
    output STAT_TX_PACKET_64_BYTES;
    output STAT_TX_PACKET_65_127_BYTES;
    output STAT_TX_PACKET_8192_9215_BYTES;
    output STAT_TX_PACKET_LARGE;
    output STAT_TX_PACKET_SMALL;
    output STAT_TX_PAUSE;
    output [8:0] STAT_TX_PAUSE_VALID;
    output STAT_TX_PTP_FIFO_READ_ERROR;
    output STAT_TX_PTP_FIFO_WRITE_ERROR;
    output [5:0] STAT_TX_TOTAL_BYTES;
    output [13:0] STAT_TX_TOTAL_GOOD_BYTES;
    output STAT_TX_TOTAL_GOOD_PACKETS;
    output STAT_TX_TOTAL_PACKETS;
    output STAT_TX_UNICAST;
    output STAT_TX_USER_PAUSE;
    output STAT_TX_VLAN;
    output TX_OVFOUT;
    output [4:0] TX_PTP_PCSLANE_OUT;
    output [79:0] TX_PTP_TSTAMP_OUT;
    output [15:0] TX_PTP_TSTAMP_TAG_OUT;
    output TX_PTP_TSTAMP_VALID_OUT;
    output TX_RDYOUT;
    output [15:0] TX_SERDES_ALT_DATA0;
    output [15:0] TX_SERDES_ALT_DATA1;
    output [15:0] TX_SERDES_ALT_DATA2;
    output [15:0] TX_SERDES_ALT_DATA3;
    output [63:0] TX_SERDES_DATA0;
    output [63:0] TX_SERDES_DATA1;
    output [63:0] TX_SERDES_DATA2;
    output [63:0] TX_SERDES_DATA3;
    output [31:0] TX_SERDES_DATA4;
    output [31:0] TX_SERDES_DATA5;
    output [31:0] TX_SERDES_DATA6;
    output [31:0] TX_SERDES_DATA7;
    output [31:0] TX_SERDES_DATA8;
    output [31:0] TX_SERDES_DATA9;
    output TX_UNFOUT;
    input CTL_CAUI4_MODE;
    input CTL_RSFEC_ENABLE_TRANSCODER_BYPASS_MODE;
    input CTL_RSFEC_IEEE_ERROR_INDICATION_MODE;
    input CTL_RX_CHECK_ETYPE_GCP;
    input CTL_RX_CHECK_ETYPE_GPP;
    input CTL_RX_CHECK_ETYPE_PCP;
    input CTL_RX_CHECK_ETYPE_PPP;
    input CTL_RX_CHECK_MCAST_GCP;
    input CTL_RX_CHECK_MCAST_GPP;
    input CTL_RX_CHECK_MCAST_PCP;
    input CTL_RX_CHECK_MCAST_PPP;
    input CTL_RX_CHECK_OPCODE_GCP;
    input CTL_RX_CHECK_OPCODE_GPP;
    input CTL_RX_CHECK_OPCODE_PCP;
    input CTL_RX_CHECK_OPCODE_PPP;
    input CTL_RX_CHECK_SA_GCP;
    input CTL_RX_CHECK_SA_GPP;
    input CTL_RX_CHECK_SA_PCP;
    input CTL_RX_CHECK_SA_PPP;
    input CTL_RX_CHECK_UCAST_GCP;
    input CTL_RX_CHECK_UCAST_GPP;
    input CTL_RX_CHECK_UCAST_PCP;
    input CTL_RX_CHECK_UCAST_PPP;
    input CTL_RX_ENABLE;
    input CTL_RX_ENABLE_GCP;
    input CTL_RX_ENABLE_GPP;
    input CTL_RX_ENABLE_PCP;
    input CTL_RX_ENABLE_PPP;
    input CTL_RX_FORCE_RESYNC;
    input [8:0] CTL_RX_PAUSE_ACK;
    input [8:0] CTL_RX_PAUSE_ENABLE;
    input CTL_RX_RSFEC_ENABLE;
    input CTL_RX_RSFEC_ENABLE_CORRECTION;
    input CTL_RX_RSFEC_ENABLE_INDICATION;
    input [79:0] CTL_RX_SYSTEMTIMERIN;
    input CTL_RX_TEST_PATTERN;
    input CTL_TX_ENABLE;
    input CTL_TX_LANE0_VLM_BIP7_OVERRIDE;
    input [7:0] CTL_TX_LANE0_VLM_BIP7_OVERRIDE_VALUE;
    input [8:0] CTL_TX_PAUSE_ENABLE;
    input [15:0] CTL_TX_PAUSE_QUANTA0;
    input [15:0] CTL_TX_PAUSE_QUANTA1;
    input [15:0] CTL_TX_PAUSE_QUANTA2;
    input [15:0] CTL_TX_PAUSE_QUANTA3;
    input [15:0] CTL_TX_PAUSE_QUANTA4;
    input [15:0] CTL_TX_PAUSE_QUANTA5;
    input [15:0] CTL_TX_PAUSE_QUANTA6;
    input [15:0] CTL_TX_PAUSE_QUANTA7;
    input [15:0] CTL_TX_PAUSE_QUANTA8;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER0;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER1;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER2;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER3;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER4;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER5;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER6;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER7;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER8;
    input [8:0] CTL_TX_PAUSE_REQ;
    input CTL_TX_PTP_VLANE_ADJUST_MODE;
    input CTL_TX_RESEND_PAUSE;
    input CTL_TX_RSFEC_ENABLE;
    input CTL_TX_SEND_IDLE;
    input CTL_TX_SEND_LFI;
    input CTL_TX_SEND_RFI;
    input [79:0] CTL_TX_SYSTEMTIMERIN;
    input CTL_TX_TEST_PATTERN;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input [329:0] RSFEC_BYPASS_RX_DIN;
    input RSFEC_BYPASS_RX_DIN_CW_START;
    input [329:0] RSFEC_BYPASS_TX_DIN;
    input RSFEC_BYPASS_TX_DIN_CW_START;
    input RX_CLK;
    input RX_RESET;
    input [15:0] RX_SERDES_ALT_DATA0;
    input [15:0] RX_SERDES_ALT_DATA1;
    input [15:0] RX_SERDES_ALT_DATA2;
    input [15:0] RX_SERDES_ALT_DATA3;
    input [9:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA0;
    input [63:0] RX_SERDES_DATA1;
    input [63:0] RX_SERDES_DATA2;
    input [63:0] RX_SERDES_DATA3;
    input [31:0] RX_SERDES_DATA4;
    input [31:0] RX_SERDES_DATA5;
    input [31:0] RX_SERDES_DATA6;
    input [31:0] RX_SERDES_DATA7;
    input [31:0] RX_SERDES_DATA8;
    input [31:0] RX_SERDES_DATA9;
    input [9:0] RX_SERDES_RESET;
    input TX_CLK;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input [55:0] TX_PREIN;
    input [1:0] TX_PTP_1588OP_IN;
    input [15:0] TX_PTP_CHKSUM_OFFSET_IN;
    input [63:0] TX_PTP_RXTSTAMP_IN;
    input [15:0] TX_PTP_TAG_FIELD_IN;
    input [15:0] TX_PTP_TSTAMP_OFFSET_IN;
    input TX_PTP_UPD_CHKSUM_IN;
    input TX_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module PPC405_ADV (...);
    parameter in_delay=100;
    parameter out_delay=100;
    output APUFCMDECODED;
    output APUFCMDECUDIVALID;
    output APUFCMENDIAN;
    output APUFCMFLUSH;
    output APUFCMINSTRVALID;
    output APUFCMLOADDVALID;
    output APUFCMOPERANDVALID;
    output APUFCMWRITEBACKOK;
    output APUFCMXERCA;
    output C405CPMCORESLEEPREQ;
    output C405CPMMSRCE;
    output C405CPMMSREE;
    output C405CPMTIMERIRQ;
    output C405CPMTIMERRESETREQ;
    output C405DBGLOADDATAONAPUDBUS;
    output C405DBGMSRWE;
    output C405DBGSTOPACK;
    output C405DBGWBCOMPLETE;
    output C405DBGWBFULL;
    output C405JTGCAPTUREDR;
    output C405JTGEXTEST;
    output C405JTGPGMOUT;
    output C405JTGSHIFTDR;
    output C405JTGTDO;
    output C405JTGTDOEN;
    output C405JTGUPDATEDR;
    output C405PLBDCUABORT;
    output C405PLBDCUCACHEABLE;
    output C405PLBDCUGUARDED;
    output C405PLBDCUREQUEST;
    output C405PLBDCURNW;
    output C405PLBDCUSIZE2;
    output C405PLBDCUU0ATTR;
    output C405PLBDCUWRITETHRU;
    output C405PLBICUABORT;
    output C405PLBICUCACHEABLE;
    output C405PLBICUREQUEST;
    output C405PLBICUU0ATTR;
    output C405RSTCHIPRESETREQ;
    output C405RSTCORERESETREQ;
    output C405RSTSYSRESETREQ;
    output C405TRCCYCLE;
    output C405TRCTRIGGEREVENTOUT;
    output C405XXXMACHINECHECK;
    output DCREMACCLK;
    output DCREMACENABLER;
    output DCREMACREAD;
    output DCREMACWRITE;
    output DSOCMBRAMEN;
    output DSOCMBUSY;
    output DSOCMRDADDRVALID;
    output DSOCMWRADDRVALID;
    output EXTDCRREAD;
    output EXTDCRWRITE;
    output ISOCMBRAMEN;
    output ISOCMBRAMEVENWRITEEN;
    output ISOCMBRAMODDWRITEEN;
    output ISOCMDCRBRAMEVENEN;
    output ISOCMDCRBRAMODDEN;
    output ISOCMDCRBRAMRDSELECT;
    output [0:10] C405TRCTRIGGEREVENTTYPE;
    output [0:1] C405PLBDCUPRIORITY;
    output [0:1] C405PLBICUPRIORITY;
    output [0:1] C405TRCEVENEXECUTIONSTATUS;
    output [0:1] C405TRCODDEXECUTIONSTATUS;
    output [0:29] C405DBGWBIAR;
    output [0:29] C405PLBICUABUS;
    output [0:2] APUFCMDECUDI;
    output [0:31] APUFCMINSTRUCTION;
    output [0:31] APUFCMLOADDATA;
    output [0:31] APUFCMRADATA;
    output [0:31] APUFCMRBDATA;
    output [0:31] C405PLBDCUABUS;
    output [0:31] DCREMACDBUS;
    output [0:31] DSOCMBRAMWRDBUS;
    output [0:31] EXTDCRDBUSOUT;
    output [0:31] ISOCMBRAMWRDBUS;
    output [0:3] APUFCMLOADBYTEEN;
    output [0:3] C405TRCTRACESTATUS;
    output [0:3] DSOCMBRAMBYTEWRITE;
    output [0:63] C405PLBDCUWRDBUS;
    output [0:7] C405PLBDCUBE;
    output [0:9] EXTDCRABUS;
    output [2:3] C405PLBICUSIZE;
    output [8:28] ISOCMBRAMRDABUS;
    output [8:28] ISOCMBRAMWRABUS;
    output [8:29] DSOCMBRAMABUS;
    output [8:9] DCREMACABUS;
    input BRAMDSOCMCLK;
    input BRAMISOCMCLK;
    input CPMC405CLOCK;
    input CPMC405CORECLKINACTIVE;
    input CPMC405CPUCLKEN;
    input CPMC405JTAGCLKEN;
    input CPMC405SYNCBYPASS;
    input CPMC405TIMERCLKEN;
    input CPMC405TIMERTICK;
    input CPMDCRCLK;
    input CPMFCMCLK;
    input DBGC405DEBUGHALT;
    input DBGC405EXTBUSHOLDACK;
    input DBGC405UNCONDDEBUGEVENT;
    input DSOCMRWCOMPLETE;
    input EICC405CRITINPUTIRQ;
    input EICC405EXTINPUTIRQ;
    input EMACDCRACK;
    input EXTDCRACK;
    input FCMAPUDCDCREN;
    input FCMAPUDCDFORCEALIGN;
    input FCMAPUDCDFORCEBESTEERING;
    input FCMAPUDCDFPUOP;
    input FCMAPUDCDGPRWRITE;
    input FCMAPUDCDLDSTBYTE;
    input FCMAPUDCDLDSTDW;
    input FCMAPUDCDLDSTHW;
    input FCMAPUDCDLDSTQW;
    input FCMAPUDCDLDSTWD;
    input FCMAPUDCDLOAD;
    input FCMAPUDCDPRIVOP;
    input FCMAPUDCDRAEN;
    input FCMAPUDCDRBEN;
    input FCMAPUDCDSTORE;
    input FCMAPUDCDTRAPBE;
    input FCMAPUDCDTRAPLE;
    input FCMAPUDCDUPDATE;
    input FCMAPUDCDXERCAEN;
    input FCMAPUDCDXEROVEN;
    input FCMAPUDECODEBUSY;
    input FCMAPUDONE;
    input FCMAPUEXCEPTION;
    input FCMAPUEXEBLOCKINGMCO;
    input FCMAPUEXENONBLOCKINGMCO;
    input FCMAPUINSTRACK;
    input FCMAPULOADWAIT;
    input FCMAPURESULTVALID;
    input FCMAPUSLEEPNOTREADY;
    input FCMAPUXERCA;
    input FCMAPUXEROV;
    input JTGC405BNDSCANTDO;
    input JTGC405TCK;
    input JTGC405TDI;
    input JTGC405TMS;
    input JTGC405TRSTNEG;
    input MCBCPUCLKEN;
    input MCBJTAGEN;
    input MCBTIMEREN;
    input MCPPCRST;
    input PLBC405DCUADDRACK;
    input PLBC405DCUBUSY;
    input PLBC405DCUERR;
    input PLBC405DCURDDACK;
    input PLBC405DCUSSIZE1;
    input PLBC405DCUWRDACK;
    input PLBC405ICUADDRACK;
    input PLBC405ICUBUSY;
    input PLBC405ICUERR;
    input PLBC405ICURDDACK;
    input PLBC405ICUSSIZE1;
    input PLBCLK;
    input RSTC405RESETCHIP;
    input RSTC405RESETCORE;
    input RSTC405RESETSYS;
    input TIEC405DETERMINISTICMULT;
    input TIEC405DISOPERANDFWD;
    input TIEC405MMUEN;
    input TIEPVRBIT10;
    input TIEPVRBIT11;
    input TIEPVRBIT28;
    input TIEPVRBIT29;
    input TIEPVRBIT30;
    input TIEPVRBIT31;
    input TIEPVRBIT8;
    input TIEPVRBIT9;
    input TRCC405TRACEDISABLE;
    input TRCC405TRIGGEREVENTIN;
    input [0:15] TIEAPUCONTROL;
    input [0:23] TIEAPUUDI1;
    input [0:23] TIEAPUUDI2;
    input [0:23] TIEAPUUDI3;
    input [0:23] TIEAPUUDI4;
    input [0:23] TIEAPUUDI5;
    input [0:23] TIEAPUUDI6;
    input [0:23] TIEAPUUDI7;
    input [0:23] TIEAPUUDI8;
    input [0:2] FCMAPUEXECRFIELD;
    input [0:31] BRAMDSOCMRDDBUS;
    input [0:31] BRAMISOCMDCRRDDBUS;
    input [0:31] EMACDCRDBUS;
    input [0:31] EXTDCRDBUSIN;
    input [0:31] FCMAPURESULT;
    input [0:3] FCMAPUCR;
    input [0:5] TIEDCRADDR;
    input [0:63] BRAMISOCMRDDBUS;
    input [0:63] PLBC405DCURDDBUS;
    input [0:63] PLBC405ICURDDBUS;
    input [0:7] DSARCVALUE;
    input [0:7] DSCNTLVALUE;
    input [0:7] ISARCVALUE;
    input [0:7] ISCNTLVALUE;
    input [1:3] PLBC405DCURDWDADDR;
    input [1:3] PLBC405ICURDWDADDR;
endmodule

module PPC440 (...);
    parameter CLOCK_DELAY = "FALSE";
    parameter DCR_AUTOLOCK_ENABLE = "TRUE";
    parameter PPCDM_ASYNCMODE = "FALSE";
    parameter PPCDS_ASYNCMODE = "FALSE";
    parameter PPCS0_WIDTH_128N64 = "TRUE";
    parameter PPCS1_WIDTH_128N64 = "TRUE";
    parameter [0:16] APU_CONTROL = 17'h02000;
    parameter [0:23] APU_UDI0 = 24'h000000;
    parameter [0:23] APU_UDI1 = 24'h000000;
    parameter [0:23] APU_UDI10 = 24'h000000;
    parameter [0:23] APU_UDI11 = 24'h000000;
    parameter [0:23] APU_UDI12 = 24'h000000;
    parameter [0:23] APU_UDI13 = 24'h000000;
    parameter [0:23] APU_UDI14 = 24'h000000;
    parameter [0:23] APU_UDI15 = 24'h000000;
    parameter [0:23] APU_UDI2 = 24'h000000;
    parameter [0:23] APU_UDI3 = 24'h000000;
    parameter [0:23] APU_UDI4 = 24'h000000;
    parameter [0:23] APU_UDI5 = 24'h000000;
    parameter [0:23] APU_UDI6 = 24'h000000;
    parameter [0:23] APU_UDI7 = 24'h000000;
    parameter [0:23] APU_UDI8 = 24'h000000;
    parameter [0:23] APU_UDI9 = 24'h000000;
    parameter [0:31] DMA0_RXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA0_TXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA1_RXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA1_TXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA2_RXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA2_TXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA3_RXCHANNELCTRL = 32'h01010000;
    parameter [0:31] DMA3_TXCHANNELCTRL = 32'h01010000;
    parameter [0:31] INTERCONNECT_IMASK = 32'hFFFFFFFF;
    parameter [0:31] INTERCONNECT_TMPL_SEL = 32'h3FFFFFFF;
    parameter [0:31] MI_ARBCONFIG = 32'h00432010;
    parameter [0:31] MI_BANKCONFLICT_MASK = 32'h00000000;
    parameter [0:31] MI_CONTROL = 32'h0000008F;
    parameter [0:31] MI_ROWCONFLICT_MASK = 32'h00000000;
    parameter [0:31] PPCM_ARBCONFIG = 32'h00432010;
    parameter [0:31] PPCM_CONTROL = 32'h8000019F;
    parameter [0:31] PPCM_COUNTER = 32'h00000500;
    parameter [0:31] PPCS0_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
    parameter [0:31] PPCS0_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
    parameter [0:31] PPCS0_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
    parameter [0:31] PPCS0_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
    parameter [0:31] PPCS0_CONTROL = 32'h8033336C;
    parameter [0:31] PPCS1_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
    parameter [0:31] PPCS1_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
    parameter [0:31] PPCS1_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
    parameter [0:31] PPCS1_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
    parameter [0:31] PPCS1_CONTROL = 32'h8033336C;
    parameter [0:31] XBAR_ADDRMAP_TMPL0 = 32'hFFFF0000;
    parameter [0:31] XBAR_ADDRMAP_TMPL1 = 32'h00000000;
    parameter [0:31] XBAR_ADDRMAP_TMPL2 = 32'h00000000;
    parameter [0:31] XBAR_ADDRMAP_TMPL3 = 32'h00000000;
    parameter [0:7] DMA0_CONTROL = 8'h00;
    parameter [0:7] DMA1_CONTROL = 8'h00;
    parameter [0:7] DMA2_CONTROL = 8'h00;
    parameter [0:7] DMA3_CONTROL = 8'h00;
    parameter [0:9] DMA0_RXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA0_TXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA1_RXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA1_TXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA2_RXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA2_TXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA3_RXIRQTIMER = 10'h3FF;
    parameter [0:9] DMA3_TXIRQTIMER = 10'h3FF;
    output APUFCMDECFPUOP;
    output APUFCMDECLOAD;
    output APUFCMDECNONAUTON;
    output APUFCMDECSTORE;
    output APUFCMDECUDIVALID;
    output APUFCMENDIAN;
    output APUFCMFLUSH;
    output APUFCMINSTRVALID;
    output APUFCMLOADDVALID;
    output APUFCMMSRFE0;
    output APUFCMMSRFE1;
    output APUFCMNEXTINSTRREADY;
    output APUFCMOPERANDVALID;
    output APUFCMWRITEBACKOK;
    output C440CPMCORESLEEPREQ;
    output C440CPMDECIRPTREQ;
    output C440CPMFITIRPTREQ;
    output C440CPMMSRCE;
    output C440CPMMSREE;
    output C440CPMTIMERRESETREQ;
    output C440CPMWDIRPTREQ;
    output C440JTGTDO;
    output C440JTGTDOEN;
    output C440MACHINECHECK;
    output C440RSTCHIPRESETREQ;
    output C440RSTCORERESETREQ;
    output C440RSTSYSTEMRESETREQ;
    output C440TRCCYCLE;
    output C440TRCTRIGGEREVENTOUT;
    output DMA0LLRSTENGINEACK;
    output DMA0LLRXDSTRDYN;
    output DMA0LLTXEOFN;
    output DMA0LLTXEOPN;
    output DMA0LLTXSOFN;
    output DMA0LLTXSOPN;
    output DMA0LLTXSRCRDYN;
    output DMA0RXIRQ;
    output DMA0TXIRQ;
    output DMA1LLRSTENGINEACK;
    output DMA1LLRXDSTRDYN;
    output DMA1LLTXEOFN;
    output DMA1LLTXEOPN;
    output DMA1LLTXSOFN;
    output DMA1LLTXSOPN;
    output DMA1LLTXSRCRDYN;
    output DMA1RXIRQ;
    output DMA1TXIRQ;
    output DMA2LLRSTENGINEACK;
    output DMA2LLRXDSTRDYN;
    output DMA2LLTXEOFN;
    output DMA2LLTXEOPN;
    output DMA2LLTXSOFN;
    output DMA2LLTXSOPN;
    output DMA2LLTXSRCRDYN;
    output DMA2RXIRQ;
    output DMA2TXIRQ;
    output DMA3LLRSTENGINEACK;
    output DMA3LLRXDSTRDYN;
    output DMA3LLTXEOFN;
    output DMA3LLTXEOPN;
    output DMA3LLTXSOFN;
    output DMA3LLTXSOPN;
    output DMA3LLTXSRCRDYN;
    output DMA3RXIRQ;
    output DMA3TXIRQ;
    output MIMCADDRESSVALID;
    output MIMCBANKCONFLICT;
    output MIMCREADNOTWRITE;
    output MIMCROWCONFLICT;
    output MIMCWRITEDATAVALID;
    output PPCCPMINTERCONNECTBUSY;
    output PPCDMDCRREAD;
    output PPCDMDCRWRITE;
    output PPCDSDCRACK;
    output PPCDSDCRTIMEOUTWAIT;
    output PPCEICINTERCONNECTIRQ;
    output PPCMPLBABORT;
    output PPCMPLBBUSLOCK;
    output PPCMPLBLOCKERR;
    output PPCMPLBRDBURST;
    output PPCMPLBREQUEST;
    output PPCMPLBRNW;
    output PPCMPLBWRBURST;
    output PPCS0PLBADDRACK;
    output PPCS0PLBRDBTERM;
    output PPCS0PLBRDCOMP;
    output PPCS0PLBRDDACK;
    output PPCS0PLBREARBITRATE;
    output PPCS0PLBWAIT;
    output PPCS0PLBWRBTERM;
    output PPCS0PLBWRCOMP;
    output PPCS0PLBWRDACK;
    output PPCS1PLBADDRACK;
    output PPCS1PLBRDBTERM;
    output PPCS1PLBRDCOMP;
    output PPCS1PLBRDDACK;
    output PPCS1PLBREARBITRATE;
    output PPCS1PLBWAIT;
    output PPCS1PLBWRBTERM;
    output PPCS1PLBWRCOMP;
    output PPCS1PLBWRDACK;
    output [0:127] APUFCMLOADDATA;
    output [0:127] MIMCWRITEDATA;
    output [0:127] PPCMPLBWRDBUS;
    output [0:127] PPCS0PLBRDDBUS;
    output [0:127] PPCS1PLBRDDBUS;
    output [0:13] C440TRCTRIGGEREVENTTYPE;
    output [0:15] MIMCBYTEENABLE;
    output [0:15] PPCMPLBBE;
    output [0:15] PPCMPLBTATTRIBUTE;
    output [0:1] PPCMPLBPRIORITY;
    output [0:1] PPCS0PLBSSIZE;
    output [0:1] PPCS1PLBSSIZE;
    output [0:2] APUFCMDECLDSTXFERSIZE;
    output [0:2] C440TRCBRANCHSTATUS;
    output [0:2] PPCMPLBTYPE;
    output [0:31] APUFCMINSTRUCTION;
    output [0:31] APUFCMRADATA;
    output [0:31] APUFCMRBDATA;
    output [0:31] DMA0LLTXD;
    output [0:31] DMA1LLTXD;
    output [0:31] DMA2LLTXD;
    output [0:31] DMA3LLTXD;
    output [0:31] PPCDMDCRDBUSOUT;
    output [0:31] PPCDSDCRDBUSIN;
    output [0:31] PPCMPLBABUS;
    output [0:35] MIMCADDRESS;
    output [0:3] APUFCMDECUDI;
    output [0:3] APUFCMLOADBYTEADDR;
    output [0:3] DMA0LLTXREM;
    output [0:3] DMA1LLTXREM;
    output [0:3] DMA2LLTXREM;
    output [0:3] DMA3LLTXREM;
    output [0:3] PPCMPLBSIZE;
    output [0:3] PPCS0PLBMBUSY;
    output [0:3] PPCS0PLBMIRQ;
    output [0:3] PPCS0PLBMRDERR;
    output [0:3] PPCS0PLBMWRERR;
    output [0:3] PPCS0PLBRDWDADDR;
    output [0:3] PPCS1PLBMBUSY;
    output [0:3] PPCS1PLBMIRQ;
    output [0:3] PPCS1PLBMRDERR;
    output [0:3] PPCS1PLBMWRERR;
    output [0:3] PPCS1PLBRDWDADDR;
    output [0:4] C440TRCEXECUTIONSTATUS;
    output [0:6] C440TRCTRACESTATUS;
    output [0:7] C440DBGSYSTEMCONTROL;
    output [0:9] PPCDMDCRABUS;
    output [20:21] PPCDMDCRUABUS;
    output [28:31] PPCMPLBUABUS;
    input CPMC440CLK;
    input CPMC440CLKEN;
    input CPMC440CORECLOCKINACTIVE;
    input CPMC440TIMERCLOCK;
    input CPMDCRCLK;
    input CPMDMA0LLCLK;
    input CPMDMA1LLCLK;
    input CPMDMA2LLCLK;
    input CPMDMA3LLCLK;
    input CPMFCMCLK;
    input CPMINTERCONNECTCLK;
    input CPMINTERCONNECTCLKEN;
    input CPMINTERCONNECTCLKNTO1;
    input CPMMCCLK;
    input CPMPPCMPLBCLK;
    input CPMPPCS0PLBCLK;
    input CPMPPCS1PLBCLK;
    input DBGC440DEBUGHALT;
    input DBGC440UNCONDDEBUGEVENT;
    input DCRPPCDMACK;
    input DCRPPCDMTIMEOUTWAIT;
    input DCRPPCDSREAD;
    input DCRPPCDSWRITE;
    input EICC440CRITIRQ;
    input EICC440EXTIRQ;
    input FCMAPUCONFIRMINSTR;
    input FCMAPUDONE;
    input FCMAPUEXCEPTION;
    input FCMAPUFPSCRFEX;
    input FCMAPURESULTVALID;
    input FCMAPUSLEEPNOTREADY;
    input JTGC440TCK;
    input JTGC440TDI;
    input JTGC440TMS;
    input JTGC440TRSTNEG;
    input LLDMA0RSTENGINEREQ;
    input LLDMA0RXEOFN;
    input LLDMA0RXEOPN;
    input LLDMA0RXSOFN;
    input LLDMA0RXSOPN;
    input LLDMA0RXSRCRDYN;
    input LLDMA0TXDSTRDYN;
    input LLDMA1RSTENGINEREQ;
    input LLDMA1RXEOFN;
    input LLDMA1RXEOPN;
    input LLDMA1RXSOFN;
    input LLDMA1RXSOPN;
    input LLDMA1RXSRCRDYN;
    input LLDMA1TXDSTRDYN;
    input LLDMA2RSTENGINEREQ;
    input LLDMA2RXEOFN;
    input LLDMA2RXEOPN;
    input LLDMA2RXSOFN;
    input LLDMA2RXSOPN;
    input LLDMA2RXSRCRDYN;
    input LLDMA2TXDSTRDYN;
    input LLDMA3RSTENGINEREQ;
    input LLDMA3RXEOFN;
    input LLDMA3RXEOPN;
    input LLDMA3RXSOFN;
    input LLDMA3RXSOPN;
    input LLDMA3RXSRCRDYN;
    input LLDMA3TXDSTRDYN;
    input MCMIADDRREADYTOACCEPT;
    input MCMIREADDATAERR;
    input MCMIREADDATAVALID;
    input PLBPPCMADDRACK;
    input PLBPPCMMBUSY;
    input PLBPPCMMIRQ;
    input PLBPPCMMRDERR;
    input PLBPPCMMWRERR;
    input PLBPPCMRDBTERM;
    input PLBPPCMRDDACK;
    input PLBPPCMRDPENDREQ;
    input PLBPPCMREARBITRATE;
    input PLBPPCMTIMEOUT;
    input PLBPPCMWRBTERM;
    input PLBPPCMWRDACK;
    input PLBPPCMWRPENDREQ;
    input PLBPPCS0ABORT;
    input PLBPPCS0BUSLOCK;
    input PLBPPCS0LOCKERR;
    input PLBPPCS0PAVALID;
    input PLBPPCS0RDBURST;
    input PLBPPCS0RDPENDREQ;
    input PLBPPCS0RDPRIM;
    input PLBPPCS0RNW;
    input PLBPPCS0SAVALID;
    input PLBPPCS0WRBURST;
    input PLBPPCS0WRPENDREQ;
    input PLBPPCS0WRPRIM;
    input PLBPPCS1ABORT;
    input PLBPPCS1BUSLOCK;
    input PLBPPCS1LOCKERR;
    input PLBPPCS1PAVALID;
    input PLBPPCS1RDBURST;
    input PLBPPCS1RDPENDREQ;
    input PLBPPCS1RDPRIM;
    input PLBPPCS1RNW;
    input PLBPPCS1SAVALID;
    input PLBPPCS1WRBURST;
    input PLBPPCS1WRPENDREQ;
    input PLBPPCS1WRPRIM;
    input RSTC440RESETCHIP;
    input RSTC440RESETCORE;
    input RSTC440RESETSYSTEM;
    input TIEC440ENDIANRESET;
    input TRCC440TRACEDISABLE;
    input TRCC440TRIGGEREVENTIN;
    input [0:127] FCMAPUSTOREDATA;
    input [0:127] MCMIREADDATA;
    input [0:127] PLBPPCMRDDBUS;
    input [0:127] PLBPPCS0WRDBUS;
    input [0:127] PLBPPCS1WRDBUS;
    input [0:15] PLBPPCS0BE;
    input [0:15] PLBPPCS0TATTRIBUTE;
    input [0:15] PLBPPCS1BE;
    input [0:15] PLBPPCS1TATTRIBUTE;
    input [0:1] PLBPPCMRDPENDPRI;
    input [0:1] PLBPPCMREQPRI;
    input [0:1] PLBPPCMSSIZE;
    input [0:1] PLBPPCMWRPENDPRI;
    input [0:1] PLBPPCS0MASTERID;
    input [0:1] PLBPPCS0MSIZE;
    input [0:1] PLBPPCS0RDPENDPRI;
    input [0:1] PLBPPCS0REQPRI;
    input [0:1] PLBPPCS0WRPENDPRI;
    input [0:1] PLBPPCS1MASTERID;
    input [0:1] PLBPPCS1MSIZE;
    input [0:1] PLBPPCS1RDPENDPRI;
    input [0:1] PLBPPCS1REQPRI;
    input [0:1] PLBPPCS1WRPENDPRI;
    input [0:1] TIEC440DCURDLDCACHEPLBPRIO;
    input [0:1] TIEC440DCURDNONCACHEPLBPRIO;
    input [0:1] TIEC440DCURDTOUCHPLBPRIO;
    input [0:1] TIEC440DCURDURGENTPLBPRIO;
    input [0:1] TIEC440DCUWRFLUSHPLBPRIO;
    input [0:1] TIEC440DCUWRSTOREPLBPRIO;
    input [0:1] TIEC440DCUWRURGENTPLBPRIO;
    input [0:1] TIEC440ICURDFETCHPLBPRIO;
    input [0:1] TIEC440ICURDSPECPLBPRIO;
    input [0:1] TIEC440ICURDTOUCHPLBPRIO;
    input [0:1] TIEDCRBASEADDR;
    input [0:2] PLBPPCS0TYPE;
    input [0:2] PLBPPCS1TYPE;
    input [0:31] DCRPPCDMDBUSIN;
    input [0:31] DCRPPCDSDBUSOUT;
    input [0:31] FCMAPURESULT;
    input [0:31] LLDMA0RXD;
    input [0:31] LLDMA1RXD;
    input [0:31] LLDMA2RXD;
    input [0:31] LLDMA3RXD;
    input [0:31] PLBPPCS0ABUS;
    input [0:31] PLBPPCS1ABUS;
    input [0:3] FCMAPUCR;
    input [0:3] LLDMA0RXREM;
    input [0:3] LLDMA1RXREM;
    input [0:3] LLDMA2RXREM;
    input [0:3] LLDMA3RXREM;
    input [0:3] PLBPPCMRDWDADDR;
    input [0:3] PLBPPCS0SIZE;
    input [0:3] PLBPPCS1SIZE;
    input [0:3] TIEC440ERPNRESET;
    input [0:3] TIEC440USERRESET;
    input [0:4] DBGC440SYSTEMSTATUS;
    input [0:9] DCRPPCDSABUS;
    input [28:31] PLBPPCS0UABUS;
    input [28:31] PLBPPCS1UABUS;
    input [28:31] TIEC440PIR;
    input [28:31] TIEC440PVR;
endmodule

module MCB (...);
    parameter integer ARB_NUM_TIME_SLOTS = 12;
    parameter [17:0] ARB_TIME_SLOT_0 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_1 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_10 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_11 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_2 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_3 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_4 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_5 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_6 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_7 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_8 = 18'b111111111111111111;
    parameter [17:0] ARB_TIME_SLOT_9 = 18'b111111111111111111;
    parameter [2:0] CAL_BA = 3'h0;
    parameter CAL_BYPASS = "YES";
    parameter [11:0] CAL_CA = 12'h000;
    parameter CAL_CALIBRATION_MODE = "NOCALIBRATION";
    parameter integer CAL_CLK_DIV = 1;
    parameter CAL_DELAY = "QUARTER";
    parameter [14:0] CAL_RA = 15'h0000;
    parameter MEM_ADDR_ORDER = "BANK_ROW_COLUMN";
    parameter integer MEM_BA_SIZE = 3;
    parameter integer MEM_BURST_LEN = 8;
    parameter integer MEM_CAS_LATENCY = 4;
    parameter integer MEM_CA_SIZE = 11;
    parameter MEM_DDR1_2_ODS = "FULL";
    parameter MEM_DDR2_3_HIGH_TEMP_SR = "NORMAL";
    parameter MEM_DDR2_3_PA_SR = "FULL";
    parameter integer MEM_DDR2_ADD_LATENCY = 0;
    parameter MEM_DDR2_DIFF_DQS_EN = "YES";
    parameter MEM_DDR2_RTT = "50OHMS";
    parameter integer MEM_DDR2_WRT_RECOVERY = 4;
    parameter MEM_DDR3_ADD_LATENCY = "OFF";
    parameter MEM_DDR3_AUTO_SR = "ENABLED";
    parameter integer MEM_DDR3_CAS_LATENCY = 7;
    parameter integer MEM_DDR3_CAS_WR_LATENCY = 5;
    parameter MEM_DDR3_DYN_WRT_ODT = "OFF";
    parameter MEM_DDR3_ODS = "DIV7";
    parameter MEM_DDR3_RTT = "DIV2";
    parameter integer MEM_DDR3_WRT_RECOVERY = 7;
    parameter MEM_MDDR_ODS = "FULL";
    parameter MEM_MOBILE_PA_SR = "FULL";
    parameter integer MEM_MOBILE_TC_SR = 0;
    parameter integer MEM_RAS_VAL = 0;
    parameter integer MEM_RA_SIZE = 13;
    parameter integer MEM_RCD_VAL = 1;
    parameter integer MEM_REFI_VAL = 0;
    parameter integer MEM_RFC_VAL = 0;
    parameter integer MEM_RP_VAL = 0;
    parameter integer MEM_RTP_VAL = 0;
    parameter MEM_TYPE = "DDR3";
    parameter integer MEM_WIDTH = 4;
    parameter integer MEM_WR_VAL = 0;
    parameter integer MEM_WTR_VAL = 3;
    parameter PORT_CONFIG = "B32_B32_B32_B32";
    output CAS;
    output CKE;
    output DQIOWEN0;
    output DQSIOWEN90N;
    output DQSIOWEN90P;
    output IOIDRPADD;
    output IOIDRPBROADCAST;
    output IOIDRPCLK;
    output IOIDRPCS;
    output IOIDRPSDO;
    output IOIDRPTRAIN;
    output IOIDRPUPDATE;
    output LDMN;
    output LDMP;
    output ODT;
    output P0CMDEMPTY;
    output P0CMDFULL;
    output P0RDEMPTY;
    output P0RDERROR;
    output P0RDFULL;
    output P0RDOVERFLOW;
    output P0WREMPTY;
    output P0WRERROR;
    output P0WRFULL;
    output P0WRUNDERRUN;
    output P1CMDEMPTY;
    output P1CMDFULL;
    output P1RDEMPTY;
    output P1RDERROR;
    output P1RDFULL;
    output P1RDOVERFLOW;
    output P1WREMPTY;
    output P1WRERROR;
    output P1WRFULL;
    output P1WRUNDERRUN;
    output P2CMDEMPTY;
    output P2CMDFULL;
    output P2EMPTY;
    output P2ERROR;
    output P2FULL;
    output P2RDOVERFLOW;
    output P2WRUNDERRUN;
    output P3CMDEMPTY;
    output P3CMDFULL;
    output P3EMPTY;
    output P3ERROR;
    output P3FULL;
    output P3RDOVERFLOW;
    output P3WRUNDERRUN;
    output P4CMDEMPTY;
    output P4CMDFULL;
    output P4EMPTY;
    output P4ERROR;
    output P4FULL;
    output P4RDOVERFLOW;
    output P4WRUNDERRUN;
    output P5CMDEMPTY;
    output P5CMDFULL;
    output P5EMPTY;
    output P5ERROR;
    output P5FULL;
    output P5RDOVERFLOW;
    output P5WRUNDERRUN;
    output RAS;
    output RST;
    output SELFREFRESHMODE;
    output UDMN;
    output UDMP;
    output UOCALSTART;
    output UOCMDREADYIN;
    output UODATAVALID;
    output UODONECAL;
    output UOREFRSHFLAG;
    output UOSDO;
    output WE;
    output [14:0] ADDR;
    output [15:0] DQON;
    output [15:0] DQOP;
    output [2:0] BA;
    output [31:0] P0RDDATA;
    output [31:0] P1RDDATA;
    output [31:0] P2RDDATA;
    output [31:0] P3RDDATA;
    output [31:0] P4RDDATA;
    output [31:0] P5RDDATA;
    output [31:0] STATUS;
    output [4:0] IOIDRPADDR;
    output [6:0] P0RDCOUNT;
    output [6:0] P0WRCOUNT;
    output [6:0] P1RDCOUNT;
    output [6:0] P1WRCOUNT;
    output [6:0] P2COUNT;
    output [6:0] P3COUNT;
    output [6:0] P4COUNT;
    output [6:0] P5COUNT;
    output [7:0] UODATA;
    input DQSIOIN;
    input DQSIOIP;
    input IOIDRPSDI;
    input P0ARBEN;
    input P0CMDCLK;
    input P0CMDEN;
    input P0RDCLK;
    input P0RDEN;
    input P0WRCLK;
    input P0WREN;
    input P1ARBEN;
    input P1CMDCLK;
    input P1CMDEN;
    input P1RDCLK;
    input P1RDEN;
    input P1WRCLK;
    input P1WREN;
    input P2ARBEN;
    input P2CLK;
    input P2CMDCLK;
    input P2CMDEN;
    input P2EN;
    input P3ARBEN;
    input P3CLK;
    input P3CMDCLK;
    input P3CMDEN;
    input P3EN;
    input P4ARBEN;
    input P4CLK;
    input P4CMDCLK;
    input P4CMDEN;
    input P4EN;
    input P5ARBEN;
    input P5CLK;
    input P5CMDCLK;
    input P5CMDEN;
    input P5EN;
    input PLLLOCK;
    input RECAL;
    input SELFREFRESHENTER;
    input SYSRST;
    input UDQSIOIN;
    input UDQSIOIP;
    input UIADD;
    input UIBROADCAST;
    input UICLK;
    input UICMD;
    input UICMDEN;
    input UICMDIN;
    input UICS;
    input UIDONECAL;
    input UIDQLOWERDEC;
    input UIDQLOWERINC;
    input UIDQUPPERDEC;
    input UIDQUPPERINC;
    input UIDRPUPDATE;
    input UILDQSDEC;
    input UILDQSINC;
    input UIREAD;
    input UISDI;
    input UIUDQSDEC;
    input UIUDQSINC;
    input [11:0] P0CMDCA;
    input [11:0] P1CMDCA;
    input [11:0] P2CMDCA;
    input [11:0] P3CMDCA;
    input [11:0] P4CMDCA;
    input [11:0] P5CMDCA;
    input [14:0] P0CMDRA;
    input [14:0] P1CMDRA;
    input [14:0] P2CMDRA;
    input [14:0] P3CMDRA;
    input [14:0] P4CMDRA;
    input [14:0] P5CMDRA;
    input [15:0] DQI;
    input [1:0] PLLCE;
    input [1:0] PLLCLK;
    input [2:0] P0CMDBA;
    input [2:0] P0CMDINSTR;
    input [2:0] P1CMDBA;
    input [2:0] P1CMDINSTR;
    input [2:0] P2CMDBA;
    input [2:0] P2CMDINSTR;
    input [2:0] P3CMDBA;
    input [2:0] P3CMDINSTR;
    input [2:0] P4CMDBA;
    input [2:0] P4CMDINSTR;
    input [2:0] P5CMDBA;
    input [2:0] P5CMDINSTR;
    input [31:0] P0WRDATA;
    input [31:0] P1WRDATA;
    input [31:0] P2WRDATA;
    input [31:0] P3WRDATA;
    input [31:0] P4WRDATA;
    input [31:0] P5WRDATA;
    input [3:0] P0RWRMASK;
    input [3:0] P1RWRMASK;
    input [3:0] P2WRMASK;
    input [3:0] P3WRMASK;
    input [3:0] P4WRMASK;
    input [3:0] P5WRMASK;
    input [3:0] UIDQCOUNT;
    input [4:0] UIADDR;
    input [5:0] P0CMDBL;
    input [5:0] P1CMDBL;
    input [5:0] P2CMDBL;
    input [5:0] P3CMDBL;
    input [5:0] P4CMDBL;
    input [5:0] P5CMDBL;
endmodule

(* keep *)
module PS7 (...);
    output DMA0DAVALID;
    output DMA0DRREADY;
    output DMA0RSTN;
    output DMA1DAVALID;
    output DMA1DRREADY;
    output DMA1RSTN;
    output DMA2DAVALID;
    output DMA2DRREADY;
    output DMA2RSTN;
    output DMA3DAVALID;
    output DMA3DRREADY;
    output DMA3RSTN;
    output EMIOCAN0PHYTX;
    output EMIOCAN1PHYTX;
    output EMIOENET0GMIITXEN;
    output EMIOENET0GMIITXER;
    output EMIOENET0MDIOMDC;
    output EMIOENET0MDIOO;
    output EMIOENET0MDIOTN;
    output EMIOENET0PTPDELAYREQRX;
    output EMIOENET0PTPDELAYREQTX;
    output EMIOENET0PTPPDELAYREQRX;
    output EMIOENET0PTPPDELAYREQTX;
    output EMIOENET0PTPPDELAYRESPRX;
    output EMIOENET0PTPPDELAYRESPTX;
    output EMIOENET0PTPSYNCFRAMERX;
    output EMIOENET0PTPSYNCFRAMETX;
    output EMIOENET0SOFRX;
    output EMIOENET0SOFTX;
    output EMIOENET1GMIITXEN;
    output EMIOENET1GMIITXER;
    output EMIOENET1MDIOMDC;
    output EMIOENET1MDIOO;
    output EMIOENET1MDIOTN;
    output EMIOENET1PTPDELAYREQRX;
    output EMIOENET1PTPDELAYREQTX;
    output EMIOENET1PTPPDELAYREQRX;
    output EMIOENET1PTPPDELAYREQTX;
    output EMIOENET1PTPPDELAYRESPRX;
    output EMIOENET1PTPPDELAYRESPTX;
    output EMIOENET1PTPSYNCFRAMERX;
    output EMIOENET1PTPSYNCFRAMETX;
    output EMIOENET1SOFRX;
    output EMIOENET1SOFTX;
    output EMIOI2C0SCLO;
    output EMIOI2C0SCLTN;
    output EMIOI2C0SDAO;
    output EMIOI2C0SDATN;
    output EMIOI2C1SCLO;
    output EMIOI2C1SCLTN;
    output EMIOI2C1SDAO;
    output EMIOI2C1SDATN;
    output EMIOPJTAGTDO;
    output EMIOPJTAGTDTN;
    output EMIOSDIO0BUSPOW;
    output EMIOSDIO0CLK;
    output EMIOSDIO0CMDO;
    output EMIOSDIO0CMDTN;
    output EMIOSDIO0LED;
    output EMIOSDIO1BUSPOW;
    output EMIOSDIO1CLK;
    output EMIOSDIO1CMDO;
    output EMIOSDIO1CMDTN;
    output EMIOSDIO1LED;
    output EMIOSPI0MO;
    output EMIOSPI0MOTN;
    output EMIOSPI0SCLKO;
    output EMIOSPI0SCLKTN;
    output EMIOSPI0SO;
    output EMIOSPI0SSNTN;
    output EMIOSPI0STN;
    output EMIOSPI1MO;
    output EMIOSPI1MOTN;
    output EMIOSPI1SCLKO;
    output EMIOSPI1SCLKTN;
    output EMIOSPI1SO;
    output EMIOSPI1SSNTN;
    output EMIOSPI1STN;
    output EMIOTRACECTL;
    output EMIOUART0DTRN;
    output EMIOUART0RTSN;
    output EMIOUART0TX;
    output EMIOUART1DTRN;
    output EMIOUART1RTSN;
    output EMIOUART1TX;
    output EMIOUSB0VBUSPWRSELECT;
    output EMIOUSB1VBUSPWRSELECT;
    output EMIOWDTRSTO;
    output EVENTEVENTO;
    output MAXIGP0ARESETN;
    output MAXIGP0ARVALID;
    output MAXIGP0AWVALID;
    output MAXIGP0BREADY;
    output MAXIGP0RREADY;
    output MAXIGP0WLAST;
    output MAXIGP0WVALID;
    output MAXIGP1ARESETN;
    output MAXIGP1ARVALID;
    output MAXIGP1AWVALID;
    output MAXIGP1BREADY;
    output MAXIGP1RREADY;
    output MAXIGP1WLAST;
    output MAXIGP1WVALID;
    output SAXIACPARESETN;
    output SAXIACPARREADY;
    output SAXIACPAWREADY;
    output SAXIACPBVALID;
    output SAXIACPRLAST;
    output SAXIACPRVALID;
    output SAXIACPWREADY;
    output SAXIGP0ARESETN;
    output SAXIGP0ARREADY;
    output SAXIGP0AWREADY;
    output SAXIGP0BVALID;
    output SAXIGP0RLAST;
    output SAXIGP0RVALID;
    output SAXIGP0WREADY;
    output SAXIGP1ARESETN;
    output SAXIGP1ARREADY;
    output SAXIGP1AWREADY;
    output SAXIGP1BVALID;
    output SAXIGP1RLAST;
    output SAXIGP1RVALID;
    output SAXIGP1WREADY;
    output SAXIHP0ARESETN;
    output SAXIHP0ARREADY;
    output SAXIHP0AWREADY;
    output SAXIHP0BVALID;
    output SAXIHP0RLAST;
    output SAXIHP0RVALID;
    output SAXIHP0WREADY;
    output SAXIHP1ARESETN;
    output SAXIHP1ARREADY;
    output SAXIHP1AWREADY;
    output SAXIHP1BVALID;
    output SAXIHP1RLAST;
    output SAXIHP1RVALID;
    output SAXIHP1WREADY;
    output SAXIHP2ARESETN;
    output SAXIHP2ARREADY;
    output SAXIHP2AWREADY;
    output SAXIHP2BVALID;
    output SAXIHP2RLAST;
    output SAXIHP2RVALID;
    output SAXIHP2WREADY;
    output SAXIHP3ARESETN;
    output SAXIHP3ARREADY;
    output SAXIHP3AWREADY;
    output SAXIHP3BVALID;
    output SAXIHP3RLAST;
    output SAXIHP3RVALID;
    output SAXIHP3WREADY;
    output [11:0] MAXIGP0ARID;
    output [11:0] MAXIGP0AWID;
    output [11:0] MAXIGP0WID;
    output [11:0] MAXIGP1ARID;
    output [11:0] MAXIGP1AWID;
    output [11:0] MAXIGP1WID;
    output [1:0] DMA0DATYPE;
    output [1:0] DMA1DATYPE;
    output [1:0] DMA2DATYPE;
    output [1:0] DMA3DATYPE;
    output [1:0] EMIOUSB0PORTINDCTL;
    output [1:0] EMIOUSB1PORTINDCTL;
    output [1:0] EVENTSTANDBYWFE;
    output [1:0] EVENTSTANDBYWFI;
    output [1:0] MAXIGP0ARBURST;
    output [1:0] MAXIGP0ARLOCK;
    output [1:0] MAXIGP0ARSIZE;
    output [1:0] MAXIGP0AWBURST;
    output [1:0] MAXIGP0AWLOCK;
    output [1:0] MAXIGP0AWSIZE;
    output [1:0] MAXIGP1ARBURST;
    output [1:0] MAXIGP1ARLOCK;
    output [1:0] MAXIGP1ARSIZE;
    output [1:0] MAXIGP1AWBURST;
    output [1:0] MAXIGP1AWLOCK;
    output [1:0] MAXIGP1AWSIZE;
    output [1:0] SAXIACPBRESP;
    output [1:0] SAXIACPRRESP;
    output [1:0] SAXIGP0BRESP;
    output [1:0] SAXIGP0RRESP;
    output [1:0] SAXIGP1BRESP;
    output [1:0] SAXIGP1RRESP;
    output [1:0] SAXIHP0BRESP;
    output [1:0] SAXIHP0RRESP;
    output [1:0] SAXIHP1BRESP;
    output [1:0] SAXIHP1RRESP;
    output [1:0] SAXIHP2BRESP;
    output [1:0] SAXIHP2RRESP;
    output [1:0] SAXIHP3BRESP;
    output [1:0] SAXIHP3RRESP;
    output [28:0] IRQP2F;
    output [2:0] EMIOSDIO0BUSVOLT;
    output [2:0] EMIOSDIO1BUSVOLT;
    output [2:0] EMIOSPI0SSON;
    output [2:0] EMIOSPI1SSON;
    output [2:0] EMIOTTC0WAVEO;
    output [2:0] EMIOTTC1WAVEO;
    output [2:0] MAXIGP0ARPROT;
    output [2:0] MAXIGP0AWPROT;
    output [2:0] MAXIGP1ARPROT;
    output [2:0] MAXIGP1AWPROT;
    output [2:0] SAXIACPBID;
    output [2:0] SAXIACPRID;
    output [2:0] SAXIHP0RACOUNT;
    output [2:0] SAXIHP1RACOUNT;
    output [2:0] SAXIHP2RACOUNT;
    output [2:0] SAXIHP3RACOUNT;
    output [31:0] EMIOTRACEDATA;
    output [31:0] FTMTP2FDEBUG;
    output [31:0] MAXIGP0ARADDR;
    output [31:0] MAXIGP0AWADDR;
    output [31:0] MAXIGP0WDATA;
    output [31:0] MAXIGP1ARADDR;
    output [31:0] MAXIGP1AWADDR;
    output [31:0] MAXIGP1WDATA;
    output [31:0] SAXIGP0RDATA;
    output [31:0] SAXIGP1RDATA;
    output [3:0] EMIOSDIO0DATAO;
    output [3:0] EMIOSDIO0DATATN;
    output [3:0] EMIOSDIO1DATAO;
    output [3:0] EMIOSDIO1DATATN;
    output [3:0] FCLKCLK;
    output [3:0] FCLKRESETN;
    output [3:0] FTMTF2PTRIGACK;
    output [3:0] FTMTP2FTRIG;
    output [3:0] MAXIGP0ARCACHE;
    output [3:0] MAXIGP0ARLEN;
    output [3:0] MAXIGP0ARQOS;
    output [3:0] MAXIGP0AWCACHE;
    output [3:0] MAXIGP0AWLEN;
    output [3:0] MAXIGP0AWQOS;
    output [3:0] MAXIGP0WSTRB;
    output [3:0] MAXIGP1ARCACHE;
    output [3:0] MAXIGP1ARLEN;
    output [3:0] MAXIGP1ARQOS;
    output [3:0] MAXIGP1AWCACHE;
    output [3:0] MAXIGP1AWLEN;
    output [3:0] MAXIGP1AWQOS;
    output [3:0] MAXIGP1WSTRB;
    output [5:0] SAXIGP0BID;
    output [5:0] SAXIGP0RID;
    output [5:0] SAXIGP1BID;
    output [5:0] SAXIGP1RID;
    output [5:0] SAXIHP0BID;
    output [5:0] SAXIHP0RID;
    output [5:0] SAXIHP0WACOUNT;
    output [5:0] SAXIHP1BID;
    output [5:0] SAXIHP1RID;
    output [5:0] SAXIHP1WACOUNT;
    output [5:0] SAXIHP2BID;
    output [5:0] SAXIHP2RID;
    output [5:0] SAXIHP2WACOUNT;
    output [5:0] SAXIHP3BID;
    output [5:0] SAXIHP3RID;
    output [5:0] SAXIHP3WACOUNT;
    output [63:0] EMIOGPIOO;
    output [63:0] EMIOGPIOTN;
    output [63:0] SAXIACPRDATA;
    output [63:0] SAXIHP0RDATA;
    output [63:0] SAXIHP1RDATA;
    output [63:0] SAXIHP2RDATA;
    output [63:0] SAXIHP3RDATA;
    output [7:0] EMIOENET0GMIITXD;
    output [7:0] EMIOENET1GMIITXD;
    output [7:0] SAXIHP0RCOUNT;
    output [7:0] SAXIHP0WCOUNT;
    output [7:0] SAXIHP1RCOUNT;
    output [7:0] SAXIHP1WCOUNT;
    output [7:0] SAXIHP2RCOUNT;
    output [7:0] SAXIHP2WCOUNT;
    output [7:0] SAXIHP3RCOUNT;
    output [7:0] SAXIHP3WCOUNT;
    inout DDRCASB;
    inout DDRCKE;
    inout DDRCKN;
    inout DDRCKP;
    inout DDRCSB;
    inout DDRDRSTB;
    inout DDRODT;
    inout DDRRASB;
    inout DDRVRN;
    inout DDRVRP;
    inout DDRWEB;
    inout PSCLK;
    inout PSPORB;
    inout PSSRSTB;
    inout [14:0] DDRA;
    inout [2:0] DDRBA;
    inout [31:0] DDRDQ;
    inout [3:0] DDRDM;
    inout [3:0] DDRDQSN;
    inout [3:0] DDRDQSP;
    inout [53:0] MIO;
    input DMA0ACLK;
    input DMA0DAREADY;
    input DMA0DRLAST;
    input DMA0DRVALID;
    input DMA1ACLK;
    input DMA1DAREADY;
    input DMA1DRLAST;
    input DMA1DRVALID;
    input DMA2ACLK;
    input DMA2DAREADY;
    input DMA2DRLAST;
    input DMA2DRVALID;
    input DMA3ACLK;
    input DMA3DAREADY;
    input DMA3DRLAST;
    input DMA3DRVALID;
    input EMIOCAN0PHYRX;
    input EMIOCAN1PHYRX;
    input EMIOENET0EXTINTIN;
    input EMIOENET0GMIICOL;
    input EMIOENET0GMIICRS;
    input EMIOENET0GMIIRXCLK;
    input EMIOENET0GMIIRXDV;
    input EMIOENET0GMIIRXER;
    input EMIOENET0GMIITXCLK;
    input EMIOENET0MDIOI;
    input EMIOENET1EXTINTIN;
    input EMIOENET1GMIICOL;
    input EMIOENET1GMIICRS;
    input EMIOENET1GMIIRXCLK;
    input EMIOENET1GMIIRXDV;
    input EMIOENET1GMIIRXER;
    input EMIOENET1GMIITXCLK;
    input EMIOENET1MDIOI;
    input EMIOI2C0SCLI;
    input EMIOI2C0SDAI;
    input EMIOI2C1SCLI;
    input EMIOI2C1SDAI;
    input EMIOPJTAGTCK;
    input EMIOPJTAGTDI;
    input EMIOPJTAGTMS;
    input EMIOSDIO0CDN;
    input EMIOSDIO0CLKFB;
    input EMIOSDIO0CMDI;
    input EMIOSDIO0WP;
    input EMIOSDIO1CDN;
    input EMIOSDIO1CLKFB;
    input EMIOSDIO1CMDI;
    input EMIOSDIO1WP;
    input EMIOSPI0MI;
    input EMIOSPI0SCLKI;
    input EMIOSPI0SI;
    input EMIOSPI0SSIN;
    input EMIOSPI1MI;
    input EMIOSPI1SCLKI;
    input EMIOSPI1SI;
    input EMIOSPI1SSIN;
    input EMIOSRAMINTIN;
    input EMIOTRACECLK;
    input EMIOUART0CTSN;
    input EMIOUART0DCDN;
    input EMIOUART0DSRN;
    input EMIOUART0RIN;
    input EMIOUART0RX;
    input EMIOUART1CTSN;
    input EMIOUART1DCDN;
    input EMIOUART1DSRN;
    input EMIOUART1RIN;
    input EMIOUART1RX;
    input EMIOUSB0VBUSPWRFAULT;
    input EMIOUSB1VBUSPWRFAULT;
    input EMIOWDTCLKI;
    input EVENTEVENTI;
    input FPGAIDLEN;
    input FTMDTRACEINCLOCK;
    input FTMDTRACEINVALID;
    input MAXIGP0ACLK;
    input MAXIGP0ARREADY;
    input MAXIGP0AWREADY;
    input MAXIGP0BVALID;
    input MAXIGP0RLAST;
    input MAXIGP0RVALID;
    input MAXIGP0WREADY;
    input MAXIGP1ACLK;
    input MAXIGP1ARREADY;
    input MAXIGP1AWREADY;
    input MAXIGP1BVALID;
    input MAXIGP1RLAST;
    input MAXIGP1RVALID;
    input MAXIGP1WREADY;
    input SAXIACPACLK;
    input SAXIACPARVALID;
    input SAXIACPAWVALID;
    input SAXIACPBREADY;
    input SAXIACPRREADY;
    input SAXIACPWLAST;
    input SAXIACPWVALID;
    input SAXIGP0ACLK;
    input SAXIGP0ARVALID;
    input SAXIGP0AWVALID;
    input SAXIGP0BREADY;
    input SAXIGP0RREADY;
    input SAXIGP0WLAST;
    input SAXIGP0WVALID;
    input SAXIGP1ACLK;
    input SAXIGP1ARVALID;
    input SAXIGP1AWVALID;
    input SAXIGP1BREADY;
    input SAXIGP1RREADY;
    input SAXIGP1WLAST;
    input SAXIGP1WVALID;
    input SAXIHP0ACLK;
    input SAXIHP0ARVALID;
    input SAXIHP0AWVALID;
    input SAXIHP0BREADY;
    input SAXIHP0RDISSUECAP1EN;
    input SAXIHP0RREADY;
    input SAXIHP0WLAST;
    input SAXIHP0WRISSUECAP1EN;
    input SAXIHP0WVALID;
    input SAXIHP1ACLK;
    input SAXIHP1ARVALID;
    input SAXIHP1AWVALID;
    input SAXIHP1BREADY;
    input SAXIHP1RDISSUECAP1EN;
    input SAXIHP1RREADY;
    input SAXIHP1WLAST;
    input SAXIHP1WRISSUECAP1EN;
    input SAXIHP1WVALID;
    input SAXIHP2ACLK;
    input SAXIHP2ARVALID;
    input SAXIHP2AWVALID;
    input SAXIHP2BREADY;
    input SAXIHP2RDISSUECAP1EN;
    input SAXIHP2RREADY;
    input SAXIHP2WLAST;
    input SAXIHP2WRISSUECAP1EN;
    input SAXIHP2WVALID;
    input SAXIHP3ACLK;
    input SAXIHP3ARVALID;
    input SAXIHP3AWVALID;
    input SAXIHP3BREADY;
    input SAXIHP3RDISSUECAP1EN;
    input SAXIHP3RREADY;
    input SAXIHP3WLAST;
    input SAXIHP3WRISSUECAP1EN;
    input SAXIHP3WVALID;
    input [11:0] MAXIGP0BID;
    input [11:0] MAXIGP0RID;
    input [11:0] MAXIGP1BID;
    input [11:0] MAXIGP1RID;
    input [19:0] IRQF2P;
    input [1:0] DMA0DRTYPE;
    input [1:0] DMA1DRTYPE;
    input [1:0] DMA2DRTYPE;
    input [1:0] DMA3DRTYPE;
    input [1:0] MAXIGP0BRESP;
    input [1:0] MAXIGP0RRESP;
    input [1:0] MAXIGP1BRESP;
    input [1:0] MAXIGP1RRESP;
    input [1:0] SAXIACPARBURST;
    input [1:0] SAXIACPARLOCK;
    input [1:0] SAXIACPARSIZE;
    input [1:0] SAXIACPAWBURST;
    input [1:0] SAXIACPAWLOCK;
    input [1:0] SAXIACPAWSIZE;
    input [1:0] SAXIGP0ARBURST;
    input [1:0] SAXIGP0ARLOCK;
    input [1:0] SAXIGP0ARSIZE;
    input [1:0] SAXIGP0AWBURST;
    input [1:0] SAXIGP0AWLOCK;
    input [1:0] SAXIGP0AWSIZE;
    input [1:0] SAXIGP1ARBURST;
    input [1:0] SAXIGP1ARLOCK;
    input [1:0] SAXIGP1ARSIZE;
    input [1:0] SAXIGP1AWBURST;
    input [1:0] SAXIGP1AWLOCK;
    input [1:0] SAXIGP1AWSIZE;
    input [1:0] SAXIHP0ARBURST;
    input [1:0] SAXIHP0ARLOCK;
    input [1:0] SAXIHP0ARSIZE;
    input [1:0] SAXIHP0AWBURST;
    input [1:0] SAXIHP0AWLOCK;
    input [1:0] SAXIHP0AWSIZE;
    input [1:0] SAXIHP1ARBURST;
    input [1:0] SAXIHP1ARLOCK;
    input [1:0] SAXIHP1ARSIZE;
    input [1:0] SAXIHP1AWBURST;
    input [1:0] SAXIHP1AWLOCK;
    input [1:0] SAXIHP1AWSIZE;
    input [1:0] SAXIHP2ARBURST;
    input [1:0] SAXIHP2ARLOCK;
    input [1:0] SAXIHP2ARSIZE;
    input [1:0] SAXIHP2AWBURST;
    input [1:0] SAXIHP2AWLOCK;
    input [1:0] SAXIHP2AWSIZE;
    input [1:0] SAXIHP3ARBURST;
    input [1:0] SAXIHP3ARLOCK;
    input [1:0] SAXIHP3ARSIZE;
    input [1:0] SAXIHP3AWBURST;
    input [1:0] SAXIHP3AWLOCK;
    input [1:0] SAXIHP3AWSIZE;
    input [2:0] EMIOTTC0CLKI;
    input [2:0] EMIOTTC1CLKI;
    input [2:0] SAXIACPARID;
    input [2:0] SAXIACPARPROT;
    input [2:0] SAXIACPAWID;
    input [2:0] SAXIACPAWPROT;
    input [2:0] SAXIACPWID;
    input [2:0] SAXIGP0ARPROT;
    input [2:0] SAXIGP0AWPROT;
    input [2:0] SAXIGP1ARPROT;
    input [2:0] SAXIGP1AWPROT;
    input [2:0] SAXIHP0ARPROT;
    input [2:0] SAXIHP0AWPROT;
    input [2:0] SAXIHP1ARPROT;
    input [2:0] SAXIHP1AWPROT;
    input [2:0] SAXIHP2ARPROT;
    input [2:0] SAXIHP2AWPROT;
    input [2:0] SAXIHP3ARPROT;
    input [2:0] SAXIHP3AWPROT;
    input [31:0] FTMDTRACEINDATA;
    input [31:0] FTMTF2PDEBUG;
    input [31:0] MAXIGP0RDATA;
    input [31:0] MAXIGP1RDATA;
    input [31:0] SAXIACPARADDR;
    input [31:0] SAXIACPAWADDR;
    input [31:0] SAXIGP0ARADDR;
    input [31:0] SAXIGP0AWADDR;
    input [31:0] SAXIGP0WDATA;
    input [31:0] SAXIGP1ARADDR;
    input [31:0] SAXIGP1AWADDR;
    input [31:0] SAXIGP1WDATA;
    input [31:0] SAXIHP0ARADDR;
    input [31:0] SAXIHP0AWADDR;
    input [31:0] SAXIHP1ARADDR;
    input [31:0] SAXIHP1AWADDR;
    input [31:0] SAXIHP2ARADDR;
    input [31:0] SAXIHP2AWADDR;
    input [31:0] SAXIHP3ARADDR;
    input [31:0] SAXIHP3AWADDR;
    input [3:0] DDRARB;
    input [3:0] EMIOSDIO0DATAI;
    input [3:0] EMIOSDIO1DATAI;
    input [3:0] FCLKCLKTRIGN;
    input [3:0] FTMDTRACEINATID;
    input [3:0] FTMTF2PTRIG;
    input [3:0] FTMTP2FTRIGACK;
    input [3:0] SAXIACPARCACHE;
    input [3:0] SAXIACPARLEN;
    input [3:0] SAXIACPARQOS;
    input [3:0] SAXIACPAWCACHE;
    input [3:0] SAXIACPAWLEN;
    input [3:0] SAXIACPAWQOS;
    input [3:0] SAXIGP0ARCACHE;
    input [3:0] SAXIGP0ARLEN;
    input [3:0] SAXIGP0ARQOS;
    input [3:0] SAXIGP0AWCACHE;
    input [3:0] SAXIGP0AWLEN;
    input [3:0] SAXIGP0AWQOS;
    input [3:0] SAXIGP0WSTRB;
    input [3:0] SAXIGP1ARCACHE;
    input [3:0] SAXIGP1ARLEN;
    input [3:0] SAXIGP1ARQOS;
    input [3:0] SAXIGP1AWCACHE;
    input [3:0] SAXIGP1AWLEN;
    input [3:0] SAXIGP1AWQOS;
    input [3:0] SAXIGP1WSTRB;
    input [3:0] SAXIHP0ARCACHE;
    input [3:0] SAXIHP0ARLEN;
    input [3:0] SAXIHP0ARQOS;
    input [3:0] SAXIHP0AWCACHE;
    input [3:0] SAXIHP0AWLEN;
    input [3:0] SAXIHP0AWQOS;
    input [3:0] SAXIHP1ARCACHE;
    input [3:0] SAXIHP1ARLEN;
    input [3:0] SAXIHP1ARQOS;
    input [3:0] SAXIHP1AWCACHE;
    input [3:0] SAXIHP1AWLEN;
    input [3:0] SAXIHP1AWQOS;
    input [3:0] SAXIHP2ARCACHE;
    input [3:0] SAXIHP2ARLEN;
    input [3:0] SAXIHP2ARQOS;
    input [3:0] SAXIHP2AWCACHE;
    input [3:0] SAXIHP2AWLEN;
    input [3:0] SAXIHP2AWQOS;
    input [3:0] SAXIHP3ARCACHE;
    input [3:0] SAXIHP3ARLEN;
    input [3:0] SAXIHP3ARQOS;
    input [3:0] SAXIHP3AWCACHE;
    input [3:0] SAXIHP3AWLEN;
    input [3:0] SAXIHP3AWQOS;
    input [4:0] SAXIACPARUSER;
    input [4:0] SAXIACPAWUSER;
    input [5:0] SAXIGP0ARID;
    input [5:0] SAXIGP0AWID;
    input [5:0] SAXIGP0WID;
    input [5:0] SAXIGP1ARID;
    input [5:0] SAXIGP1AWID;
    input [5:0] SAXIGP1WID;
    input [5:0] SAXIHP0ARID;
    input [5:0] SAXIHP0AWID;
    input [5:0] SAXIHP0WID;
    input [5:0] SAXIHP1ARID;
    input [5:0] SAXIHP1AWID;
    input [5:0] SAXIHP1WID;
    input [5:0] SAXIHP2ARID;
    input [5:0] SAXIHP2AWID;
    input [5:0] SAXIHP2WID;
    input [5:0] SAXIHP3ARID;
    input [5:0] SAXIHP3AWID;
    input [5:0] SAXIHP3WID;
    input [63:0] EMIOGPIOI;
    input [63:0] SAXIACPWDATA;
    input [63:0] SAXIHP0WDATA;
    input [63:0] SAXIHP1WDATA;
    input [63:0] SAXIHP2WDATA;
    input [63:0] SAXIHP3WDATA;
    input [7:0] EMIOENET0GMIIRXD;
    input [7:0] EMIOENET1GMIIRXD;
    input [7:0] SAXIACPWSTRB;
    input [7:0] SAXIHP0WSTRB;
    input [7:0] SAXIHP1WSTRB;
    input [7:0] SAXIHP2WSTRB;
    input [7:0] SAXIHP3WSTRB;
endmodule

(* keep *)
module PS8 (...);
    output [7:0] ADMA2PLCACK;
    output [7:0] ADMA2PLTVLD;
    output DPAUDIOREFCLK;
    output DPAUXDATAOEN;
    output DPAUXDATAOUT;
    output DPLIVEVIDEODEOUT;
    output [31:0] DPMAXISMIXEDAUDIOTDATA;
    output DPMAXISMIXEDAUDIOTID;
    output DPMAXISMIXEDAUDIOTVALID;
    output DPSAXISAUDIOTREADY;
    output DPVIDEOOUTHSYNC;
    output [35:0] DPVIDEOOUTPIXEL1;
    output DPVIDEOOUTVSYNC;
    output DPVIDEOREFCLK;
    output EMIOCAN0PHYTX;
    output EMIOCAN1PHYTX;
    output [1:0] EMIOENET0DMABUSWIDTH;
    output EMIOENET0DMATXENDTOG;
    output [93:0] EMIOENET0GEMTSUTIMERCNT;
    output [7:0] EMIOENET0GMIITXD;
    output EMIOENET0GMIITXEN;
    output EMIOENET0GMIITXER;
    output EMIOENET0MDIOMDC;
    output EMIOENET0MDIOO;
    output EMIOENET0MDIOTN;
    output [7:0] EMIOENET0RXWDATA;
    output EMIOENET0RXWEOP;
    output EMIOENET0RXWERR;
    output EMIOENET0RXWFLUSH;
    output EMIOENET0RXWSOP;
    output [44:0] EMIOENET0RXWSTATUS;
    output EMIOENET0RXWWR;
    output [2:0] EMIOENET0SPEEDMODE;
    output EMIOENET0TXRRD;
    output [3:0] EMIOENET0TXRSTATUS;
    output [1:0] EMIOENET1DMABUSWIDTH;
    output EMIOENET1DMATXENDTOG;
    output [7:0] EMIOENET1GMIITXD;
    output EMIOENET1GMIITXEN;
    output EMIOENET1GMIITXER;
    output EMIOENET1MDIOMDC;
    output EMIOENET1MDIOO;
    output EMIOENET1MDIOTN;
    output [7:0] EMIOENET1RXWDATA;
    output EMIOENET1RXWEOP;
    output EMIOENET1RXWERR;
    output EMIOENET1RXWFLUSH;
    output EMIOENET1RXWSOP;
    output [44:0] EMIOENET1RXWSTATUS;
    output EMIOENET1RXWWR;
    output [2:0] EMIOENET1SPEEDMODE;
    output EMIOENET1TXRRD;
    output [3:0] EMIOENET1TXRSTATUS;
    output [1:0] EMIOENET2DMABUSWIDTH;
    output EMIOENET2DMATXENDTOG;
    output [7:0] EMIOENET2GMIITXD;
    output EMIOENET2GMIITXEN;
    output EMIOENET2GMIITXER;
    output EMIOENET2MDIOMDC;
    output EMIOENET2MDIOO;
    output EMIOENET2MDIOTN;
    output [7:0] EMIOENET2RXWDATA;
    output EMIOENET2RXWEOP;
    output EMIOENET2RXWERR;
    output EMIOENET2RXWFLUSH;
    output EMIOENET2RXWSOP;
    output [44:0] EMIOENET2RXWSTATUS;
    output EMIOENET2RXWWR;
    output [2:0] EMIOENET2SPEEDMODE;
    output EMIOENET2TXRRD;
    output [3:0] EMIOENET2TXRSTATUS;
    output [1:0] EMIOENET3DMABUSWIDTH;
    output EMIOENET3DMATXENDTOG;
    output [7:0] EMIOENET3GMIITXD;
    output EMIOENET3GMIITXEN;
    output EMIOENET3GMIITXER;
    output EMIOENET3MDIOMDC;
    output EMIOENET3MDIOO;
    output EMIOENET3MDIOTN;
    output [7:0] EMIOENET3RXWDATA;
    output EMIOENET3RXWEOP;
    output EMIOENET3RXWERR;
    output EMIOENET3RXWFLUSH;
    output EMIOENET3RXWSOP;
    output [44:0] EMIOENET3RXWSTATUS;
    output EMIOENET3RXWWR;
    output [2:0] EMIOENET3SPEEDMODE;
    output EMIOENET3TXRRD;
    output [3:0] EMIOENET3TXRSTATUS;
    output EMIOGEM0DELAYREQRX;
    output EMIOGEM0DELAYREQTX;
    output EMIOGEM0PDELAYREQRX;
    output EMIOGEM0PDELAYREQTX;
    output EMIOGEM0PDELAYRESPRX;
    output EMIOGEM0PDELAYRESPTX;
    output EMIOGEM0RXSOF;
    output EMIOGEM0SYNCFRAMERX;
    output EMIOGEM0SYNCFRAMETX;
    output EMIOGEM0TSUTIMERCMPVAL;
    output EMIOGEM0TXRFIXEDLAT;
    output EMIOGEM0TXSOF;
    output EMIOGEM1DELAYREQRX;
    output EMIOGEM1DELAYREQTX;
    output EMIOGEM1PDELAYREQRX;
    output EMIOGEM1PDELAYREQTX;
    output EMIOGEM1PDELAYRESPRX;
    output EMIOGEM1PDELAYRESPTX;
    output EMIOGEM1RXSOF;
    output EMIOGEM1SYNCFRAMERX;
    output EMIOGEM1SYNCFRAMETX;
    output EMIOGEM1TSUTIMERCMPVAL;
    output EMIOGEM1TXRFIXEDLAT;
    output EMIOGEM1TXSOF;
    output EMIOGEM2DELAYREQRX;
    output EMIOGEM2DELAYREQTX;
    output EMIOGEM2PDELAYREQRX;
    output EMIOGEM2PDELAYREQTX;
    output EMIOGEM2PDELAYRESPRX;
    output EMIOGEM2PDELAYRESPTX;
    output EMIOGEM2RXSOF;
    output EMIOGEM2SYNCFRAMERX;
    output EMIOGEM2SYNCFRAMETX;
    output EMIOGEM2TSUTIMERCMPVAL;
    output EMIOGEM2TXRFIXEDLAT;
    output EMIOGEM2TXSOF;
    output EMIOGEM3DELAYREQRX;
    output EMIOGEM3DELAYREQTX;
    output EMIOGEM3PDELAYREQRX;
    output EMIOGEM3PDELAYREQTX;
    output EMIOGEM3PDELAYRESPRX;
    output EMIOGEM3PDELAYRESPTX;
    output EMIOGEM3RXSOF;
    output EMIOGEM3SYNCFRAMERX;
    output EMIOGEM3SYNCFRAMETX;
    output EMIOGEM3TSUTIMERCMPVAL;
    output EMIOGEM3TXRFIXEDLAT;
    output EMIOGEM3TXSOF;
    output [95:0] EMIOGPIOO;
    output [95:0] EMIOGPIOTN;
    output EMIOI2C0SCLO;
    output EMIOI2C0SCLTN;
    output EMIOI2C0SDAO;
    output EMIOI2C0SDATN;
    output EMIOI2C1SCLO;
    output EMIOI2C1SCLTN;
    output EMIOI2C1SDAO;
    output EMIOI2C1SDATN;
    output EMIOSDIO0BUSPOWER;
    output [2:0] EMIOSDIO0BUSVOLT;
    output EMIOSDIO0CLKOUT;
    output EMIOSDIO0CMDENA;
    output EMIOSDIO0CMDOUT;
    output [7:0] EMIOSDIO0DATAENA;
    output [7:0] EMIOSDIO0DATAOUT;
    output EMIOSDIO0LEDCONTROL;
    output EMIOSDIO1BUSPOWER;
    output [2:0] EMIOSDIO1BUSVOLT;
    output EMIOSDIO1CLKOUT;
    output EMIOSDIO1CMDENA;
    output EMIOSDIO1CMDOUT;
    output [7:0] EMIOSDIO1DATAENA;
    output [7:0] EMIOSDIO1DATAOUT;
    output EMIOSDIO1LEDCONTROL;
    output EMIOSPI0MO;
    output EMIOSPI0MOTN;
    output EMIOSPI0SCLKO;
    output EMIOSPI0SCLKTN;
    output EMIOSPI0SO;
    output EMIOSPI0SSNTN;
    output [2:0] EMIOSPI0SSON;
    output EMIOSPI0STN;
    output EMIOSPI1MO;
    output EMIOSPI1MOTN;
    output EMIOSPI1SCLKO;
    output EMIOSPI1SCLKTN;
    output EMIOSPI1SO;
    output EMIOSPI1SSNTN;
    output [2:0] EMIOSPI1SSON;
    output EMIOSPI1STN;
    output [2:0] EMIOTTC0WAVEO;
    output [2:0] EMIOTTC1WAVEO;
    output [2:0] EMIOTTC2WAVEO;
    output [2:0] EMIOTTC3WAVEO;
    output EMIOU2DSPORTVBUSCTRLUSB30;
    output EMIOU2DSPORTVBUSCTRLUSB31;
    output EMIOU3DSPORTVBUSCTRLUSB30;
    output EMIOU3DSPORTVBUSCTRLUSB31;
    output EMIOUART0DTRN;
    output EMIOUART0RTSN;
    output EMIOUART0TX;
    output EMIOUART1DTRN;
    output EMIOUART1RTSN;
    output EMIOUART1TX;
    output EMIOWDT0RSTO;
    output EMIOWDT1RSTO;
    output FMIOGEM0FIFORXCLKTOPLBUFG;
    output FMIOGEM0FIFOTXCLKTOPLBUFG;
    output FMIOGEM1FIFORXCLKTOPLBUFG;
    output FMIOGEM1FIFOTXCLKTOPLBUFG;
    output FMIOGEM2FIFORXCLKTOPLBUFG;
    output FMIOGEM2FIFOTXCLKTOPLBUFG;
    output FMIOGEM3FIFORXCLKTOPLBUFG;
    output FMIOGEM3FIFOTXCLKTOPLBUFG;
    output FMIOGEMTSUCLKTOPLBUFG;
    output [31:0] FTMGPO;
    output [7:0] GDMA2PLCACK;
    output [7:0] GDMA2PLTVLD;
    output [39:0] MAXIGP0ARADDR;
    output [1:0] MAXIGP0ARBURST;
    output [3:0] MAXIGP0ARCACHE;
    output [15:0] MAXIGP0ARID;
    output [7:0] MAXIGP0ARLEN;
    output MAXIGP0ARLOCK;
    output [2:0] MAXIGP0ARPROT;
    output [3:0] MAXIGP0ARQOS;
    output [2:0] MAXIGP0ARSIZE;
    output [15:0] MAXIGP0ARUSER;
    output MAXIGP0ARVALID;
    output [39:0] MAXIGP0AWADDR;
    output [1:0] MAXIGP0AWBURST;
    output [3:0] MAXIGP0AWCACHE;
    output [15:0] MAXIGP0AWID;
    output [7:0] MAXIGP0AWLEN;
    output MAXIGP0AWLOCK;
    output [2:0] MAXIGP0AWPROT;
    output [3:0] MAXIGP0AWQOS;
    output [2:0] MAXIGP0AWSIZE;
    output [15:0] MAXIGP0AWUSER;
    output MAXIGP0AWVALID;
    output MAXIGP0BREADY;
    output MAXIGP0RREADY;
    output [127:0] MAXIGP0WDATA;
    output MAXIGP0WLAST;
    output [15:0] MAXIGP0WSTRB;
    output MAXIGP0WVALID;
    output [39:0] MAXIGP1ARADDR;
    output [1:0] MAXIGP1ARBURST;
    output [3:0] MAXIGP1ARCACHE;
    output [15:0] MAXIGP1ARID;
    output [7:0] MAXIGP1ARLEN;
    output MAXIGP1ARLOCK;
    output [2:0] MAXIGP1ARPROT;
    output [3:0] MAXIGP1ARQOS;
    output [2:0] MAXIGP1ARSIZE;
    output [15:0] MAXIGP1ARUSER;
    output MAXIGP1ARVALID;
    output [39:0] MAXIGP1AWADDR;
    output [1:0] MAXIGP1AWBURST;
    output [3:0] MAXIGP1AWCACHE;
    output [15:0] MAXIGP1AWID;
    output [7:0] MAXIGP1AWLEN;
    output MAXIGP1AWLOCK;
    output [2:0] MAXIGP1AWPROT;
    output [3:0] MAXIGP1AWQOS;
    output [2:0] MAXIGP1AWSIZE;
    output [15:0] MAXIGP1AWUSER;
    output MAXIGP1AWVALID;
    output MAXIGP1BREADY;
    output MAXIGP1RREADY;
    output [127:0] MAXIGP1WDATA;
    output MAXIGP1WLAST;
    output [15:0] MAXIGP1WSTRB;
    output MAXIGP1WVALID;
    output [39:0] MAXIGP2ARADDR;
    output [1:0] MAXIGP2ARBURST;
    output [3:0] MAXIGP2ARCACHE;
    output [15:0] MAXIGP2ARID;
    output [7:0] MAXIGP2ARLEN;
    output MAXIGP2ARLOCK;
    output [2:0] MAXIGP2ARPROT;
    output [3:0] MAXIGP2ARQOS;
    output [2:0] MAXIGP2ARSIZE;
    output [15:0] MAXIGP2ARUSER;
    output MAXIGP2ARVALID;
    output [39:0] MAXIGP2AWADDR;
    output [1:0] MAXIGP2AWBURST;
    output [3:0] MAXIGP2AWCACHE;
    output [15:0] MAXIGP2AWID;
    output [7:0] MAXIGP2AWLEN;
    output MAXIGP2AWLOCK;
    output [2:0] MAXIGP2AWPROT;
    output [3:0] MAXIGP2AWQOS;
    output [2:0] MAXIGP2AWSIZE;
    output [15:0] MAXIGP2AWUSER;
    output MAXIGP2AWVALID;
    output MAXIGP2BREADY;
    output MAXIGP2RREADY;
    output [127:0] MAXIGP2WDATA;
    output MAXIGP2WLAST;
    output [15:0] MAXIGP2WSTRB;
    output MAXIGP2WVALID;
    output OSCRTCCLK;
    output [3:0] PLCLK;
    output PMUAIBAFIFMFPDREQ;
    output PMUAIBAFIFMLPDREQ;
    output [46:0] PMUERRORTOPL;
    output [31:0] PMUPLGPO;
    output PSPLEVENTO;
    output [63:0] PSPLIRQFPD;
    output [99:0] PSPLIRQLPD;
    output [3:0] PSPLSTANDBYWFE;
    output [3:0] PSPLSTANDBYWFI;
    output PSPLTRACECTL;
    output [31:0] PSPLTRACEDATA;
    output [3:0] PSPLTRIGACK;
    output [3:0] PSPLTRIGGER;
    output PSS_ALTO_CORE_PAD_MGTTXN0OUT;
    output PSS_ALTO_CORE_PAD_MGTTXN1OUT;
    output PSS_ALTO_CORE_PAD_MGTTXN2OUT;
    output PSS_ALTO_CORE_PAD_MGTTXN3OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP0OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP1OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP2OUT;
    output PSS_ALTO_CORE_PAD_MGTTXP3OUT;
    output PSS_ALTO_CORE_PAD_PADO;
    output RPUEVENTO0;
    output RPUEVENTO1;
    output [43:0] SACEFPDACADDR;
    output [2:0] SACEFPDACPROT;
    output [3:0] SACEFPDACSNOOP;
    output SACEFPDACVALID;
    output SACEFPDARREADY;
    output SACEFPDAWREADY;
    output [5:0] SACEFPDBID;
    output [1:0] SACEFPDBRESP;
    output SACEFPDBUSER;
    output SACEFPDBVALID;
    output SACEFPDCDREADY;
    output SACEFPDCRREADY;
    output [127:0] SACEFPDRDATA;
    output [5:0] SACEFPDRID;
    output SACEFPDRLAST;
    output [3:0] SACEFPDRRESP;
    output SACEFPDRUSER;
    output SACEFPDRVALID;
    output SACEFPDWREADY;
    output SAXIACPARREADY;
    output SAXIACPAWREADY;
    output [4:0] SAXIACPBID;
    output [1:0] SAXIACPBRESP;
    output SAXIACPBVALID;
    output [127:0] SAXIACPRDATA;
    output [4:0] SAXIACPRID;
    output SAXIACPRLAST;
    output [1:0] SAXIACPRRESP;
    output SAXIACPRVALID;
    output SAXIACPWREADY;
    output SAXIGP0ARREADY;
    output SAXIGP0AWREADY;
    output [5:0] SAXIGP0BID;
    output [1:0] SAXIGP0BRESP;
    output SAXIGP0BVALID;
    output [3:0] SAXIGP0RACOUNT;
    output [7:0] SAXIGP0RCOUNT;
    output [127:0] SAXIGP0RDATA;
    output [5:0] SAXIGP0RID;
    output SAXIGP0RLAST;
    output [1:0] SAXIGP0RRESP;
    output SAXIGP0RVALID;
    output [3:0] SAXIGP0WACOUNT;
    output [7:0] SAXIGP0WCOUNT;
    output SAXIGP0WREADY;
    output SAXIGP1ARREADY;
    output SAXIGP1AWREADY;
    output [5:0] SAXIGP1BID;
    output [1:0] SAXIGP1BRESP;
    output SAXIGP1BVALID;
    output [3:0] SAXIGP1RACOUNT;
    output [7:0] SAXIGP1RCOUNT;
    output [127:0] SAXIGP1RDATA;
    output [5:0] SAXIGP1RID;
    output SAXIGP1RLAST;
    output [1:0] SAXIGP1RRESP;
    output SAXIGP1RVALID;
    output [3:0] SAXIGP1WACOUNT;
    output [7:0] SAXIGP1WCOUNT;
    output SAXIGP1WREADY;
    output SAXIGP2ARREADY;
    output SAXIGP2AWREADY;
    output [5:0] SAXIGP2BID;
    output [1:0] SAXIGP2BRESP;
    output SAXIGP2BVALID;
    output [3:0] SAXIGP2RACOUNT;
    output [7:0] SAXIGP2RCOUNT;
    output [127:0] SAXIGP2RDATA;
    output [5:0] SAXIGP2RID;
    output SAXIGP2RLAST;
    output [1:0] SAXIGP2RRESP;
    output SAXIGP2RVALID;
    output [3:0] SAXIGP2WACOUNT;
    output [7:0] SAXIGP2WCOUNT;
    output SAXIGP2WREADY;
    output SAXIGP3ARREADY;
    output SAXIGP3AWREADY;
    output [5:0] SAXIGP3BID;
    output [1:0] SAXIGP3BRESP;
    output SAXIGP3BVALID;
    output [3:0] SAXIGP3RACOUNT;
    output [7:0] SAXIGP3RCOUNT;
    output [127:0] SAXIGP3RDATA;
    output [5:0] SAXIGP3RID;
    output SAXIGP3RLAST;
    output [1:0] SAXIGP3RRESP;
    output SAXIGP3RVALID;
    output [3:0] SAXIGP3WACOUNT;
    output [7:0] SAXIGP3WCOUNT;
    output SAXIGP3WREADY;
    output SAXIGP4ARREADY;
    output SAXIGP4AWREADY;
    output [5:0] SAXIGP4BID;
    output [1:0] SAXIGP4BRESP;
    output SAXIGP4BVALID;
    output [3:0] SAXIGP4RACOUNT;
    output [7:0] SAXIGP4RCOUNT;
    output [127:0] SAXIGP4RDATA;
    output [5:0] SAXIGP4RID;
    output SAXIGP4RLAST;
    output [1:0] SAXIGP4RRESP;
    output SAXIGP4RVALID;
    output [3:0] SAXIGP4WACOUNT;
    output [7:0] SAXIGP4WCOUNT;
    output SAXIGP4WREADY;
    output SAXIGP5ARREADY;
    output SAXIGP5AWREADY;
    output [5:0] SAXIGP5BID;
    output [1:0] SAXIGP5BRESP;
    output SAXIGP5BVALID;
    output [3:0] SAXIGP5RACOUNT;
    output [7:0] SAXIGP5RCOUNT;
    output [127:0] SAXIGP5RDATA;
    output [5:0] SAXIGP5RID;
    output SAXIGP5RLAST;
    output [1:0] SAXIGP5RRESP;
    output SAXIGP5RVALID;
    output [3:0] SAXIGP5WACOUNT;
    output [7:0] SAXIGP5WCOUNT;
    output SAXIGP5WREADY;
    output SAXIGP6ARREADY;
    output SAXIGP6AWREADY;
    output [5:0] SAXIGP6BID;
    output [1:0] SAXIGP6BRESP;
    output SAXIGP6BVALID;
    output [3:0] SAXIGP6RACOUNT;
    output [7:0] SAXIGP6RCOUNT;
    output [127:0] SAXIGP6RDATA;
    output [5:0] SAXIGP6RID;
    output SAXIGP6RLAST;
    output [1:0] SAXIGP6RRESP;
    output SAXIGP6RVALID;
    output [3:0] SAXIGP6WACOUNT;
    output [7:0] SAXIGP6WCOUNT;
    output SAXIGP6WREADY;
    inout [3:0] PSS_ALTO_CORE_PAD_BOOTMODE;
    inout PSS_ALTO_CORE_PAD_CLK;
    inout PSS_ALTO_CORE_PAD_DONEB;
    inout [17:0] PSS_ALTO_CORE_PAD_DRAMA;
    inout PSS_ALTO_CORE_PAD_DRAMACTN;
    inout PSS_ALTO_CORE_PAD_DRAMALERTN;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMBA;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMBG;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCK;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCKE;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCKN;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMCSN;
    inout [8:0] PSS_ALTO_CORE_PAD_DRAMDM;
    inout [71:0] PSS_ALTO_CORE_PAD_DRAMDQ;
    inout [8:0] PSS_ALTO_CORE_PAD_DRAMDQS;
    inout [8:0] PSS_ALTO_CORE_PAD_DRAMDQSN;
    inout [1:0] PSS_ALTO_CORE_PAD_DRAMODT;
    inout PSS_ALTO_CORE_PAD_DRAMPARITY;
    inout PSS_ALTO_CORE_PAD_DRAMRAMRSTN;
    inout PSS_ALTO_CORE_PAD_ERROROUT;
    inout PSS_ALTO_CORE_PAD_ERRORSTATUS;
    inout PSS_ALTO_CORE_PAD_INITB;
    inout PSS_ALTO_CORE_PAD_JTAGTCK;
    inout PSS_ALTO_CORE_PAD_JTAGTDI;
    inout PSS_ALTO_CORE_PAD_JTAGTDO;
    inout PSS_ALTO_CORE_PAD_JTAGTMS;
    inout [77:0] PSS_ALTO_CORE_PAD_MIO;
    inout PSS_ALTO_CORE_PAD_PORB;
    inout PSS_ALTO_CORE_PAD_PROGB;
    inout PSS_ALTO_CORE_PAD_RCALIBINOUT;
    inout PSS_ALTO_CORE_PAD_SRSTB;
    inout PSS_ALTO_CORE_PAD_ZQ;
    input [7:0] ADMAFCICLK;
    input AIBPMUAFIFMFPDACK;
    input AIBPMUAFIFMLPDACK;
    input DDRCEXTREFRESHRANK0REQ;
    input DDRCEXTREFRESHRANK1REQ;
    input DDRCREFRESHPLCLK;
    input DPAUXDATAIN;
    input DPEXTERNALCUSTOMEVENT1;
    input DPEXTERNALCUSTOMEVENT2;
    input DPEXTERNALVSYNCEVENT;
    input DPHOTPLUGDETECT;
    input [7:0] DPLIVEGFXALPHAIN;
    input [35:0] DPLIVEGFXPIXEL1IN;
    input DPLIVEVIDEOINDE;
    input DPLIVEVIDEOINHSYNC;
    input [35:0] DPLIVEVIDEOINPIXEL1;
    input DPLIVEVIDEOINVSYNC;
    input DPMAXISMIXEDAUDIOTREADY;
    input DPSAXISAUDIOCLK;
    input [31:0] DPSAXISAUDIOTDATA;
    input DPSAXISAUDIOTID;
    input DPSAXISAUDIOTVALID;
    input DPVIDEOINCLK;
    input EMIOCAN0PHYRX;
    input EMIOCAN1PHYRX;
    input EMIOENET0DMATXSTATUSTOG;
    input EMIOENET0EXTINTIN;
    input EMIOENET0GMIICOL;
    input EMIOENET0GMIICRS;
    input EMIOENET0GMIIRXCLK;
    input [7:0] EMIOENET0GMIIRXD;
    input EMIOENET0GMIIRXDV;
    input EMIOENET0GMIIRXER;
    input EMIOENET0GMIITXCLK;
    input EMIOENET0MDIOI;
    input EMIOENET0RXWOVERFLOW;
    input EMIOENET0TXRCONTROL;
    input [7:0] EMIOENET0TXRDATA;
    input EMIOENET0TXRDATARDY;
    input EMIOENET0TXREOP;
    input EMIOENET0TXRERR;
    input EMIOENET0TXRFLUSHED;
    input EMIOENET0TXRSOP;
    input EMIOENET0TXRUNDERFLOW;
    input EMIOENET0TXRVALID;
    input EMIOENET1DMATXSTATUSTOG;
    input EMIOENET1EXTINTIN;
    input EMIOENET1GMIICOL;
    input EMIOENET1GMIICRS;
    input EMIOENET1GMIIRXCLK;
    input [7:0] EMIOENET1GMIIRXD;
    input EMIOENET1GMIIRXDV;
    input EMIOENET1GMIIRXER;
    input EMIOENET1GMIITXCLK;
    input EMIOENET1MDIOI;
    input EMIOENET1RXWOVERFLOW;
    input EMIOENET1TXRCONTROL;
    input [7:0] EMIOENET1TXRDATA;
    input EMIOENET1TXRDATARDY;
    input EMIOENET1TXREOP;
    input EMIOENET1TXRERR;
    input EMIOENET1TXRFLUSHED;
    input EMIOENET1TXRSOP;
    input EMIOENET1TXRUNDERFLOW;
    input EMIOENET1TXRVALID;
    input EMIOENET2DMATXSTATUSTOG;
    input EMIOENET2EXTINTIN;
    input EMIOENET2GMIICOL;
    input EMIOENET2GMIICRS;
    input EMIOENET2GMIIRXCLK;
    input [7:0] EMIOENET2GMIIRXD;
    input EMIOENET2GMIIRXDV;
    input EMIOENET2GMIIRXER;
    input EMIOENET2GMIITXCLK;
    input EMIOENET2MDIOI;
    input EMIOENET2RXWOVERFLOW;
    input EMIOENET2TXRCONTROL;
    input [7:0] EMIOENET2TXRDATA;
    input EMIOENET2TXRDATARDY;
    input EMIOENET2TXREOP;
    input EMIOENET2TXRERR;
    input EMIOENET2TXRFLUSHED;
    input EMIOENET2TXRSOP;
    input EMIOENET2TXRUNDERFLOW;
    input EMIOENET2TXRVALID;
    input EMIOENET3DMATXSTATUSTOG;
    input EMIOENET3EXTINTIN;
    input EMIOENET3GMIICOL;
    input EMIOENET3GMIICRS;
    input EMIOENET3GMIIRXCLK;
    input [7:0] EMIOENET3GMIIRXD;
    input EMIOENET3GMIIRXDV;
    input EMIOENET3GMIIRXER;
    input EMIOENET3GMIITXCLK;
    input EMIOENET3MDIOI;
    input EMIOENET3RXWOVERFLOW;
    input EMIOENET3TXRCONTROL;
    input [7:0] EMIOENET3TXRDATA;
    input EMIOENET3TXRDATARDY;
    input EMIOENET3TXREOP;
    input EMIOENET3TXRERR;
    input EMIOENET3TXRFLUSHED;
    input EMIOENET3TXRSOP;
    input EMIOENET3TXRUNDERFLOW;
    input EMIOENET3TXRVALID;
    input EMIOENETTSUCLK;
    input [1:0] EMIOGEM0TSUINCCTRL;
    input [1:0] EMIOGEM1TSUINCCTRL;
    input [1:0] EMIOGEM2TSUINCCTRL;
    input [1:0] EMIOGEM3TSUINCCTRL;
    input [95:0] EMIOGPIOI;
    input EMIOHUBPORTOVERCRNTUSB20;
    input EMIOHUBPORTOVERCRNTUSB21;
    input EMIOHUBPORTOVERCRNTUSB30;
    input EMIOHUBPORTOVERCRNTUSB31;
    input EMIOI2C0SCLI;
    input EMIOI2C0SDAI;
    input EMIOI2C1SCLI;
    input EMIOI2C1SDAI;
    input EMIOSDIO0CDN;
    input EMIOSDIO0CMDIN;
    input [7:0] EMIOSDIO0DATAIN;
    input EMIOSDIO0FBCLKIN;
    input EMIOSDIO0WP;
    input EMIOSDIO1CDN;
    input EMIOSDIO1CMDIN;
    input [7:0] EMIOSDIO1DATAIN;
    input EMIOSDIO1FBCLKIN;
    input EMIOSDIO1WP;
    input EMIOSPI0MI;
    input EMIOSPI0SCLKI;
    input EMIOSPI0SI;
    input EMIOSPI0SSIN;
    input EMIOSPI1MI;
    input EMIOSPI1SCLKI;
    input EMIOSPI1SI;
    input EMIOSPI1SSIN;
    input [2:0] EMIOTTC0CLKI;
    input [2:0] EMIOTTC1CLKI;
    input [2:0] EMIOTTC2CLKI;
    input [2:0] EMIOTTC3CLKI;
    input EMIOUART0CTSN;
    input EMIOUART0DCDN;
    input EMIOUART0DSRN;
    input EMIOUART0RIN;
    input EMIOUART0RX;
    input EMIOUART1CTSN;
    input EMIOUART1DCDN;
    input EMIOUART1DSRN;
    input EMIOUART1RIN;
    input EMIOUART1RX;
    input EMIOWDT0CLKI;
    input EMIOWDT1CLKI;
    input FMIOGEM0FIFORXCLKFROMPL;
    input FMIOGEM0FIFOTXCLKFROMPL;
    input FMIOGEM0SIGNALDETECT;
    input FMIOGEM1FIFORXCLKFROMPL;
    input FMIOGEM1FIFOTXCLKFROMPL;
    input FMIOGEM1SIGNALDETECT;
    input FMIOGEM2FIFORXCLKFROMPL;
    input FMIOGEM2FIFOTXCLKFROMPL;
    input FMIOGEM2SIGNALDETECT;
    input FMIOGEM3FIFORXCLKFROMPL;
    input FMIOGEM3FIFOTXCLKFROMPL;
    input FMIOGEM3SIGNALDETECT;
    input FMIOGEMTSUCLKFROMPL;
    input [31:0] FTMGPI;
    input [7:0] GDMAFCICLK;
    input MAXIGP0ACLK;
    input MAXIGP0ARREADY;
    input MAXIGP0AWREADY;
    input [15:0] MAXIGP0BID;
    input [1:0] MAXIGP0BRESP;
    input MAXIGP0BVALID;
    input [127:0] MAXIGP0RDATA;
    input [15:0] MAXIGP0RID;
    input MAXIGP0RLAST;
    input [1:0] MAXIGP0RRESP;
    input MAXIGP0RVALID;
    input MAXIGP0WREADY;
    input MAXIGP1ACLK;
    input MAXIGP1ARREADY;
    input MAXIGP1AWREADY;
    input [15:0] MAXIGP1BID;
    input [1:0] MAXIGP1BRESP;
    input MAXIGP1BVALID;
    input [127:0] MAXIGP1RDATA;
    input [15:0] MAXIGP1RID;
    input MAXIGP1RLAST;
    input [1:0] MAXIGP1RRESP;
    input MAXIGP1RVALID;
    input MAXIGP1WREADY;
    input MAXIGP2ACLK;
    input MAXIGP2ARREADY;
    input MAXIGP2AWREADY;
    input [15:0] MAXIGP2BID;
    input [1:0] MAXIGP2BRESP;
    input MAXIGP2BVALID;
    input [127:0] MAXIGP2RDATA;
    input [15:0] MAXIGP2RID;
    input MAXIGP2RLAST;
    input [1:0] MAXIGP2RRESP;
    input MAXIGP2RVALID;
    input MAXIGP2WREADY;
    input NFIQ0LPDRPU;
    input NFIQ1LPDRPU;
    input NIRQ0LPDRPU;
    input NIRQ1LPDRPU;
    input [7:0] PL2ADMACVLD;
    input [7:0] PL2ADMATACK;
    input [7:0] PL2GDMACVLD;
    input [7:0] PL2GDMATACK;
    input PLACECLK;
    input PLACPINACT;
    input [3:0] PLFPGASTOP;
    input [2:0] PLLAUXREFCLKFPD;
    input [1:0] PLLAUXREFCLKLPD;
    input [31:0] PLPMUGPI;
    input [3:0] PLPSAPUGICFIQ;
    input [3:0] PLPSAPUGICIRQ;
    input PLPSEVENTI;
    input [7:0] PLPSIRQ0;
    input [7:0] PLPSIRQ1;
    input PLPSTRACECLK;
    input [3:0] PLPSTRIGACK;
    input [3:0] PLPSTRIGGER;
    input [3:0] PMUERRORFROMPL;
    input PSS_ALTO_CORE_PAD_MGTRXN0IN;
    input PSS_ALTO_CORE_PAD_MGTRXN1IN;
    input PSS_ALTO_CORE_PAD_MGTRXN2IN;
    input PSS_ALTO_CORE_PAD_MGTRXN3IN;
    input PSS_ALTO_CORE_PAD_MGTRXP0IN;
    input PSS_ALTO_CORE_PAD_MGTRXP1IN;
    input PSS_ALTO_CORE_PAD_MGTRXP2IN;
    input PSS_ALTO_CORE_PAD_MGTRXP3IN;
    input PSS_ALTO_CORE_PAD_PADI;
    input PSS_ALTO_CORE_PAD_REFN0IN;
    input PSS_ALTO_CORE_PAD_REFN1IN;
    input PSS_ALTO_CORE_PAD_REFN2IN;
    input PSS_ALTO_CORE_PAD_REFN3IN;
    input PSS_ALTO_CORE_PAD_REFP0IN;
    input PSS_ALTO_CORE_PAD_REFP1IN;
    input PSS_ALTO_CORE_PAD_REFP2IN;
    input PSS_ALTO_CORE_PAD_REFP3IN;
    input RPUEVENTI0;
    input RPUEVENTI1;
    input SACEFPDACREADY;
    input [43:0] SACEFPDARADDR;
    input [1:0] SACEFPDARBAR;
    input [1:0] SACEFPDARBURST;
    input [3:0] SACEFPDARCACHE;
    input [1:0] SACEFPDARDOMAIN;
    input [5:0] SACEFPDARID;
    input [7:0] SACEFPDARLEN;
    input SACEFPDARLOCK;
    input [2:0] SACEFPDARPROT;
    input [3:0] SACEFPDARQOS;
    input [3:0] SACEFPDARREGION;
    input [2:0] SACEFPDARSIZE;
    input [3:0] SACEFPDARSNOOP;
    input [15:0] SACEFPDARUSER;
    input SACEFPDARVALID;
    input [43:0] SACEFPDAWADDR;
    input [1:0] SACEFPDAWBAR;
    input [1:0] SACEFPDAWBURST;
    input [3:0] SACEFPDAWCACHE;
    input [1:0] SACEFPDAWDOMAIN;
    input [5:0] SACEFPDAWID;
    input [7:0] SACEFPDAWLEN;
    input SACEFPDAWLOCK;
    input [2:0] SACEFPDAWPROT;
    input [3:0] SACEFPDAWQOS;
    input [3:0] SACEFPDAWREGION;
    input [2:0] SACEFPDAWSIZE;
    input [2:0] SACEFPDAWSNOOP;
    input [15:0] SACEFPDAWUSER;
    input SACEFPDAWVALID;
    input SACEFPDBREADY;
    input [127:0] SACEFPDCDDATA;
    input SACEFPDCDLAST;
    input SACEFPDCDVALID;
    input [4:0] SACEFPDCRRESP;
    input SACEFPDCRVALID;
    input SACEFPDRACK;
    input SACEFPDRREADY;
    input SACEFPDWACK;
    input [127:0] SACEFPDWDATA;
    input SACEFPDWLAST;
    input [15:0] SACEFPDWSTRB;
    input SACEFPDWUSER;
    input SACEFPDWVALID;
    input SAXIACPACLK;
    input [39:0] SAXIACPARADDR;
    input [1:0] SAXIACPARBURST;
    input [3:0] SAXIACPARCACHE;
    input [4:0] SAXIACPARID;
    input [7:0] SAXIACPARLEN;
    input SAXIACPARLOCK;
    input [2:0] SAXIACPARPROT;
    input [3:0] SAXIACPARQOS;
    input [2:0] SAXIACPARSIZE;
    input [1:0] SAXIACPARUSER;
    input SAXIACPARVALID;
    input [39:0] SAXIACPAWADDR;
    input [1:0] SAXIACPAWBURST;
    input [3:0] SAXIACPAWCACHE;
    input [4:0] SAXIACPAWID;
    input [7:0] SAXIACPAWLEN;
    input SAXIACPAWLOCK;
    input [2:0] SAXIACPAWPROT;
    input [3:0] SAXIACPAWQOS;
    input [2:0] SAXIACPAWSIZE;
    input [1:0] SAXIACPAWUSER;
    input SAXIACPAWVALID;
    input SAXIACPBREADY;
    input SAXIACPRREADY;
    input [127:0] SAXIACPWDATA;
    input SAXIACPWLAST;
    input [15:0] SAXIACPWSTRB;
    input SAXIACPWVALID;
    input [48:0] SAXIGP0ARADDR;
    input [1:0] SAXIGP0ARBURST;
    input [3:0] SAXIGP0ARCACHE;
    input [5:0] SAXIGP0ARID;
    input [7:0] SAXIGP0ARLEN;
    input SAXIGP0ARLOCK;
    input [2:0] SAXIGP0ARPROT;
    input [3:0] SAXIGP0ARQOS;
    input [2:0] SAXIGP0ARSIZE;
    input SAXIGP0ARUSER;
    input SAXIGP0ARVALID;
    input [48:0] SAXIGP0AWADDR;
    input [1:0] SAXIGP0AWBURST;
    input [3:0] SAXIGP0AWCACHE;
    input [5:0] SAXIGP0AWID;
    input [7:0] SAXIGP0AWLEN;
    input SAXIGP0AWLOCK;
    input [2:0] SAXIGP0AWPROT;
    input [3:0] SAXIGP0AWQOS;
    input [2:0] SAXIGP0AWSIZE;
    input SAXIGP0AWUSER;
    input SAXIGP0AWVALID;
    input SAXIGP0BREADY;
    input SAXIGP0RCLK;
    input SAXIGP0RREADY;
    input SAXIGP0WCLK;
    input [127:0] SAXIGP0WDATA;
    input SAXIGP0WLAST;
    input [15:0] SAXIGP0WSTRB;
    input SAXIGP0WVALID;
    input [48:0] SAXIGP1ARADDR;
    input [1:0] SAXIGP1ARBURST;
    input [3:0] SAXIGP1ARCACHE;
    input [5:0] SAXIGP1ARID;
    input [7:0] SAXIGP1ARLEN;
    input SAXIGP1ARLOCK;
    input [2:0] SAXIGP1ARPROT;
    input [3:0] SAXIGP1ARQOS;
    input [2:0] SAXIGP1ARSIZE;
    input SAXIGP1ARUSER;
    input SAXIGP1ARVALID;
    input [48:0] SAXIGP1AWADDR;
    input [1:0] SAXIGP1AWBURST;
    input [3:0] SAXIGP1AWCACHE;
    input [5:0] SAXIGP1AWID;
    input [7:0] SAXIGP1AWLEN;
    input SAXIGP1AWLOCK;
    input [2:0] SAXIGP1AWPROT;
    input [3:0] SAXIGP1AWQOS;
    input [2:0] SAXIGP1AWSIZE;
    input SAXIGP1AWUSER;
    input SAXIGP1AWVALID;
    input SAXIGP1BREADY;
    input SAXIGP1RCLK;
    input SAXIGP1RREADY;
    input SAXIGP1WCLK;
    input [127:0] SAXIGP1WDATA;
    input SAXIGP1WLAST;
    input [15:0] SAXIGP1WSTRB;
    input SAXIGP1WVALID;
    input [48:0] SAXIGP2ARADDR;
    input [1:0] SAXIGP2ARBURST;
    input [3:0] SAXIGP2ARCACHE;
    input [5:0] SAXIGP2ARID;
    input [7:0] SAXIGP2ARLEN;
    input SAXIGP2ARLOCK;
    input [2:0] SAXIGP2ARPROT;
    input [3:0] SAXIGP2ARQOS;
    input [2:0] SAXIGP2ARSIZE;
    input SAXIGP2ARUSER;
    input SAXIGP2ARVALID;
    input [48:0] SAXIGP2AWADDR;
    input [1:0] SAXIGP2AWBURST;
    input [3:0] SAXIGP2AWCACHE;
    input [5:0] SAXIGP2AWID;
    input [7:0] SAXIGP2AWLEN;
    input SAXIGP2AWLOCK;
    input [2:0] SAXIGP2AWPROT;
    input [3:0] SAXIGP2AWQOS;
    input [2:0] SAXIGP2AWSIZE;
    input SAXIGP2AWUSER;
    input SAXIGP2AWVALID;
    input SAXIGP2BREADY;
    input SAXIGP2RCLK;
    input SAXIGP2RREADY;
    input SAXIGP2WCLK;
    input [127:0] SAXIGP2WDATA;
    input SAXIGP2WLAST;
    input [15:0] SAXIGP2WSTRB;
    input SAXIGP2WVALID;
    input [48:0] SAXIGP3ARADDR;
    input [1:0] SAXIGP3ARBURST;
    input [3:0] SAXIGP3ARCACHE;
    input [5:0] SAXIGP3ARID;
    input [7:0] SAXIGP3ARLEN;
    input SAXIGP3ARLOCK;
    input [2:0] SAXIGP3ARPROT;
    input [3:0] SAXIGP3ARQOS;
    input [2:0] SAXIGP3ARSIZE;
    input SAXIGP3ARUSER;
    input SAXIGP3ARVALID;
    input [48:0] SAXIGP3AWADDR;
    input [1:0] SAXIGP3AWBURST;
    input [3:0] SAXIGP3AWCACHE;
    input [5:0] SAXIGP3AWID;
    input [7:0] SAXIGP3AWLEN;
    input SAXIGP3AWLOCK;
    input [2:0] SAXIGP3AWPROT;
    input [3:0] SAXIGP3AWQOS;
    input [2:0] SAXIGP3AWSIZE;
    input SAXIGP3AWUSER;
    input SAXIGP3AWVALID;
    input SAXIGP3BREADY;
    input SAXIGP3RCLK;
    input SAXIGP3RREADY;
    input SAXIGP3WCLK;
    input [127:0] SAXIGP3WDATA;
    input SAXIGP3WLAST;
    input [15:0] SAXIGP3WSTRB;
    input SAXIGP3WVALID;
    input [48:0] SAXIGP4ARADDR;
    input [1:0] SAXIGP4ARBURST;
    input [3:0] SAXIGP4ARCACHE;
    input [5:0] SAXIGP4ARID;
    input [7:0] SAXIGP4ARLEN;
    input SAXIGP4ARLOCK;
    input [2:0] SAXIGP4ARPROT;
    input [3:0] SAXIGP4ARQOS;
    input [2:0] SAXIGP4ARSIZE;
    input SAXIGP4ARUSER;
    input SAXIGP4ARVALID;
    input [48:0] SAXIGP4AWADDR;
    input [1:0] SAXIGP4AWBURST;
    input [3:0] SAXIGP4AWCACHE;
    input [5:0] SAXIGP4AWID;
    input [7:0] SAXIGP4AWLEN;
    input SAXIGP4AWLOCK;
    input [2:0] SAXIGP4AWPROT;
    input [3:0] SAXIGP4AWQOS;
    input [2:0] SAXIGP4AWSIZE;
    input SAXIGP4AWUSER;
    input SAXIGP4AWVALID;
    input SAXIGP4BREADY;
    input SAXIGP4RCLK;
    input SAXIGP4RREADY;
    input SAXIGP4WCLK;
    input [127:0] SAXIGP4WDATA;
    input SAXIGP4WLAST;
    input [15:0] SAXIGP4WSTRB;
    input SAXIGP4WVALID;
    input [48:0] SAXIGP5ARADDR;
    input [1:0] SAXIGP5ARBURST;
    input [3:0] SAXIGP5ARCACHE;
    input [5:0] SAXIGP5ARID;
    input [7:0] SAXIGP5ARLEN;
    input SAXIGP5ARLOCK;
    input [2:0] SAXIGP5ARPROT;
    input [3:0] SAXIGP5ARQOS;
    input [2:0] SAXIGP5ARSIZE;
    input SAXIGP5ARUSER;
    input SAXIGP5ARVALID;
    input [48:0] SAXIGP5AWADDR;
    input [1:0] SAXIGP5AWBURST;
    input [3:0] SAXIGP5AWCACHE;
    input [5:0] SAXIGP5AWID;
    input [7:0] SAXIGP5AWLEN;
    input SAXIGP5AWLOCK;
    input [2:0] SAXIGP5AWPROT;
    input [3:0] SAXIGP5AWQOS;
    input [2:0] SAXIGP5AWSIZE;
    input SAXIGP5AWUSER;
    input SAXIGP5AWVALID;
    input SAXIGP5BREADY;
    input SAXIGP5RCLK;
    input SAXIGP5RREADY;
    input SAXIGP5WCLK;
    input [127:0] SAXIGP5WDATA;
    input SAXIGP5WLAST;
    input [15:0] SAXIGP5WSTRB;
    input SAXIGP5WVALID;
    input [48:0] SAXIGP6ARADDR;
    input [1:0] SAXIGP6ARBURST;
    input [3:0] SAXIGP6ARCACHE;
    input [5:0] SAXIGP6ARID;
    input [7:0] SAXIGP6ARLEN;
    input SAXIGP6ARLOCK;
    input [2:0] SAXIGP6ARPROT;
    input [3:0] SAXIGP6ARQOS;
    input [2:0] SAXIGP6ARSIZE;
    input SAXIGP6ARUSER;
    input SAXIGP6ARVALID;
    input [48:0] SAXIGP6AWADDR;
    input [1:0] SAXIGP6AWBURST;
    input [3:0] SAXIGP6AWCACHE;
    input [5:0] SAXIGP6AWID;
    input [7:0] SAXIGP6AWLEN;
    input SAXIGP6AWLOCK;
    input [2:0] SAXIGP6AWPROT;
    input [3:0] SAXIGP6AWQOS;
    input [2:0] SAXIGP6AWSIZE;
    input SAXIGP6AWUSER;
    input SAXIGP6AWVALID;
    input SAXIGP6BREADY;
    input SAXIGP6RCLK;
    input SAXIGP6RREADY;
    input SAXIGP6WCLK;
    input [127:0] SAXIGP6WDATA;
    input SAXIGP6WLAST;
    input [15:0] SAXIGP6WSTRB;
    input SAXIGP6WVALID;
    input [59:0] STMEVENT;
endmodule

module ILKN (...);
    parameter BYPASS = "FALSE";
    parameter [1:0] CTL_RX_BURSTMAX = 2'h3;
    parameter [1:0] CTL_RX_CHAN_EXT = 2'h0;
    parameter [3:0] CTL_RX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_RX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter CTL_RX_PACKET_MODE = "TRUE";
    parameter [2:0] CTL_RX_RETRANS_MULT = 3'h0;
    parameter [3:0] CTL_RX_RETRANS_RETRY = 4'h2;
    parameter [15:0] CTL_RX_RETRANS_TIMER1 = 16'h0000;
    parameter [15:0] CTL_RX_RETRANS_TIMER2 = 16'h0008;
    parameter [11:0] CTL_RX_RETRANS_WDOG = 12'h000;
    parameter [7:0] CTL_RX_RETRANS_WRAP_TIMER = 8'h00;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [1:0] CTL_TX_BURSTMAX = 2'h3;
    parameter [2:0] CTL_TX_BURSTSHORT = 3'h1;
    parameter [1:0] CTL_TX_CHAN_EXT = 2'h0;
    parameter CTL_TX_DISABLE_SKIPWORD = "TRUE";
    parameter [6:0] CTL_TX_FC_CALLEN = 7'h00;
    parameter [3:0] CTL_TX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_TX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter [13:0] CTL_TX_RETRANS_DEPTH = 14'h0800;
    parameter [2:0] CTL_TX_RETRANS_MULT = 3'h0;
    parameter [1:0] CTL_TX_RETRANS_RAM_BANKS = 2'h3;
    parameter MODE = "TRUE";
    parameter SIM_VERSION = "2.0";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [65:0] RX_BYPASS_DATAOUT00;
    output [65:0] RX_BYPASS_DATAOUT01;
    output [65:0] RX_BYPASS_DATAOUT02;
    output [65:0] RX_BYPASS_DATAOUT03;
    output [65:0] RX_BYPASS_DATAOUT04;
    output [65:0] RX_BYPASS_DATAOUT05;
    output [65:0] RX_BYPASS_DATAOUT06;
    output [65:0] RX_BYPASS_DATAOUT07;
    output [65:0] RX_BYPASS_DATAOUT08;
    output [65:0] RX_BYPASS_DATAOUT09;
    output [65:0] RX_BYPASS_DATAOUT10;
    output [65:0] RX_BYPASS_DATAOUT11;
    output [11:0] RX_BYPASS_ENAOUT;
    output [11:0] RX_BYPASS_IS_AVAILOUT;
    output [11:0] RX_BYPASS_IS_BADLYFRAMEDOUT;
    output [11:0] RX_BYPASS_IS_OVERFLOWOUT;
    output [11:0] RX_BYPASS_IS_SYNCEDOUT;
    output [11:0] RX_BYPASS_IS_SYNCWORDOUT;
    output [10:0] RX_CHANOUT0;
    output [10:0] RX_CHANOUT1;
    output [10:0] RX_CHANOUT2;
    output [10:0] RX_CHANOUT3;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output RX_OVFOUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [11:0] STAT_RX_BAD_TYPE_ERR;
    output STAT_RX_BURSTMAX_ERR;
    output STAT_RX_BURST_ERR;
    output STAT_RX_CRC24_ERR;
    output [11:0] STAT_RX_CRC32_ERR;
    output [11:0] STAT_RX_CRC32_VALID;
    output [11:0] STAT_RX_DESCRAM_ERR;
    output [11:0] STAT_RX_DIAGWORD_INTFSTAT;
    output [11:0] STAT_RX_DIAGWORD_LANESTAT;
    output [255:0] STAT_RX_FC_STAT;
    output [11:0] STAT_RX_FRAMING_ERR;
    output STAT_RX_MEOP_ERR;
    output [11:0] STAT_RX_MF_ERR;
    output [11:0] STAT_RX_MF_LEN_ERR;
    output [11:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MSOP_ERR;
    output [7:0] STAT_RX_MUBITS;
    output STAT_RX_MUBITS_UPDATED;
    output STAT_RX_OVERFLOW_ERR;
    output STAT_RX_RETRANS_CRC24_ERR;
    output STAT_RX_RETRANS_DISC;
    output [15:0] STAT_RX_RETRANS_LATENCY;
    output STAT_RX_RETRANS_REQ;
    output STAT_RX_RETRANS_RETRY_ERR;
    output [7:0] STAT_RX_RETRANS_SEQ;
    output STAT_RX_RETRANS_SEQ_UPDATED;
    output [2:0] STAT_RX_RETRANS_STATE;
    output [4:0] STAT_RX_RETRANS_SUBSEQ;
    output STAT_RX_RETRANS_WDOG_ERR;
    output STAT_RX_RETRANS_WRAP_ERR;
    output [11:0] STAT_RX_SYNCED;
    output [11:0] STAT_RX_SYNCED_ERR;
    output [11:0] STAT_RX_WORD_SYNC;
    output STAT_TX_BURST_ERR;
    output STAT_TX_ERRINJ_BITERR_DONE;
    output STAT_TX_OVERFLOW_ERR;
    output STAT_TX_RETRANS_BURST_ERR;
    output STAT_TX_RETRANS_BUSY;
    output STAT_TX_RETRANS_RAM_PERROUT;
    output [8:0] STAT_TX_RETRANS_RAM_RADDR;
    output STAT_TX_RETRANS_RAM_RD_B0;
    output STAT_TX_RETRANS_RAM_RD_B1;
    output STAT_TX_RETRANS_RAM_RD_B2;
    output STAT_TX_RETRANS_RAM_RD_B3;
    output [1:0] STAT_TX_RETRANS_RAM_RSEL;
    output [8:0] STAT_TX_RETRANS_RAM_WADDR;
    output [643:0] STAT_TX_RETRANS_RAM_WDATA;
    output STAT_TX_RETRANS_RAM_WE_B0;
    output STAT_TX_RETRANS_RAM_WE_B1;
    output STAT_TX_RETRANS_RAM_WE_B2;
    output STAT_TX_RETRANS_RAM_WE_B3;
    output STAT_TX_UNDERFLOW_ERR;
    output TX_OVFOUT;
    output TX_RDYOUT;
    output [63:0] TX_SERDES_DATA00;
    output [63:0] TX_SERDES_DATA01;
    output [63:0] TX_SERDES_DATA02;
    output [63:0] TX_SERDES_DATA03;
    output [63:0] TX_SERDES_DATA04;
    output [63:0] TX_SERDES_DATA05;
    output [63:0] TX_SERDES_DATA06;
    output [63:0] TX_SERDES_DATA07;
    output [63:0] TX_SERDES_DATA08;
    output [63:0] TX_SERDES_DATA09;
    output [63:0] TX_SERDES_DATA10;
    output [63:0] TX_SERDES_DATA11;
    input CORE_CLK;
    input CTL_RX_FORCE_RESYNC;
    input CTL_RX_RETRANS_ACK;
    input CTL_RX_RETRANS_ENABLE;
    input CTL_RX_RETRANS_ERRIN;
    input CTL_RX_RETRANS_FORCE_REQ;
    input CTL_RX_RETRANS_RESET;
    input CTL_RX_RETRANS_RESET_MODE;
    input CTL_TX_DIAGWORD_INTFSTAT;
    input [11:0] CTL_TX_DIAGWORD_LANESTAT;
    input CTL_TX_ENABLE;
    input CTL_TX_ERRINJ_BITERR_GO;
    input [3:0] CTL_TX_ERRINJ_BITERR_LANE;
    input [255:0] CTL_TX_FC_STAT;
    input [7:0] CTL_TX_MUBITS;
    input CTL_TX_RETRANS_ENABLE;
    input CTL_TX_RETRANS_RAM_PERRIN;
    input [643:0] CTL_TX_RETRANS_RAM_RDATA;
    input CTL_TX_RETRANS_REQ;
    input CTL_TX_RETRANS_REQ_VALID;
    input [11:0] CTL_TX_RLIM_DELTA;
    input CTL_TX_RLIM_ENABLE;
    input [7:0] CTL_TX_RLIM_INTV;
    input [11:0] CTL_TX_RLIM_MAX;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input LBUS_CLK;
    input RX_BYPASS_FORCE_REALIGNIN;
    input RX_BYPASS_RDIN;
    input RX_RESET;
    input [11:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA00;
    input [63:0] RX_SERDES_DATA01;
    input [63:0] RX_SERDES_DATA02;
    input [63:0] RX_SERDES_DATA03;
    input [63:0] RX_SERDES_DATA04;
    input [63:0] RX_SERDES_DATA05;
    input [63:0] RX_SERDES_DATA06;
    input [63:0] RX_SERDES_DATA07;
    input [63:0] RX_SERDES_DATA08;
    input [63:0] RX_SERDES_DATA09;
    input [63:0] RX_SERDES_DATA10;
    input [63:0] RX_SERDES_DATA11;
    input [11:0] RX_SERDES_RESET;
    input TX_BCTLIN0;
    input TX_BCTLIN1;
    input TX_BCTLIN2;
    input TX_BCTLIN3;
    input [11:0] TX_BYPASS_CTRLIN;
    input [63:0] TX_BYPASS_DATAIN00;
    input [63:0] TX_BYPASS_DATAIN01;
    input [63:0] TX_BYPASS_DATAIN02;
    input [63:0] TX_BYPASS_DATAIN03;
    input [63:0] TX_BYPASS_DATAIN04;
    input [63:0] TX_BYPASS_DATAIN05;
    input [63:0] TX_BYPASS_DATAIN06;
    input [63:0] TX_BYPASS_DATAIN07;
    input [63:0] TX_BYPASS_DATAIN08;
    input [63:0] TX_BYPASS_DATAIN09;
    input [63:0] TX_BYPASS_DATAIN10;
    input [63:0] TX_BYPASS_DATAIN11;
    input TX_BYPASS_ENAIN;
    input [7:0] TX_BYPASS_GEARBOX_SEQIN;
    input [3:0] TX_BYPASS_MFRAMER_STATEIN;
    input [10:0] TX_CHANIN0;
    input [10:0] TX_CHANIN1;
    input [10:0] TX_CHANIN2;
    input [10:0] TX_CHANIN3;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input TX_RESET;
    input TX_SERDES_REFCLK;
    input TX_SERDES_REFCLK_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module ILKNE4 (...);
    parameter BYPASS = "FALSE";
    parameter [1:0] CTL_RX_BURSTMAX = 2'h3;
    parameter [1:0] CTL_RX_CHAN_EXT = 2'h0;
    parameter [3:0] CTL_RX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_RX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter CTL_RX_PACKET_MODE = "FALSE";
    parameter [2:0] CTL_RX_RETRANS_MULT = 3'h0;
    parameter [3:0] CTL_RX_RETRANS_RETRY = 4'h2;
    parameter [15:0] CTL_RX_RETRANS_TIMER1 = 16'h0009;
    parameter [15:0] CTL_RX_RETRANS_TIMER2 = 16'h0000;
    parameter [11:0] CTL_RX_RETRANS_WDOG = 12'h000;
    parameter [7:0] CTL_RX_RETRANS_WRAP_TIMER = 8'h00;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [1:0] CTL_TX_BURSTMAX = 2'h3;
    parameter [2:0] CTL_TX_BURSTSHORT = 3'h1;
    parameter [1:0] CTL_TX_CHAN_EXT = 2'h0;
    parameter CTL_TX_DISABLE_SKIPWORD = "FALSE";
    parameter [3:0] CTL_TX_FC_CALLEN = 4'hF;
    parameter [3:0] CTL_TX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_TX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter [13:0] CTL_TX_RETRANS_DEPTH = 14'h0800;
    parameter [2:0] CTL_TX_RETRANS_MULT = 3'h0;
    parameter [1:0] CTL_TX_RETRANS_RAM_BANKS = 2'h3;
    parameter MODE = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [65:0] RX_BYPASS_DATAOUT00;
    output [65:0] RX_BYPASS_DATAOUT01;
    output [65:0] RX_BYPASS_DATAOUT02;
    output [65:0] RX_BYPASS_DATAOUT03;
    output [65:0] RX_BYPASS_DATAOUT04;
    output [65:0] RX_BYPASS_DATAOUT05;
    output [65:0] RX_BYPASS_DATAOUT06;
    output [65:0] RX_BYPASS_DATAOUT07;
    output [65:0] RX_BYPASS_DATAOUT08;
    output [65:0] RX_BYPASS_DATAOUT09;
    output [65:0] RX_BYPASS_DATAOUT10;
    output [65:0] RX_BYPASS_DATAOUT11;
    output [11:0] RX_BYPASS_ENAOUT;
    output [11:0] RX_BYPASS_IS_AVAILOUT;
    output [11:0] RX_BYPASS_IS_BADLYFRAMEDOUT;
    output [11:0] RX_BYPASS_IS_OVERFLOWOUT;
    output [11:0] RX_BYPASS_IS_SYNCEDOUT;
    output [11:0] RX_BYPASS_IS_SYNCWORDOUT;
    output [10:0] RX_CHANOUT0;
    output [10:0] RX_CHANOUT1;
    output [10:0] RX_CHANOUT2;
    output [10:0] RX_CHANOUT3;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output RX_OVFOUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [11:0] STAT_RX_BAD_TYPE_ERR;
    output STAT_RX_BURSTMAX_ERR;
    output STAT_RX_BURST_ERR;
    output STAT_RX_CRC24_ERR;
    output [11:0] STAT_RX_CRC32_ERR;
    output [11:0] STAT_RX_CRC32_VALID;
    output [11:0] STAT_RX_DESCRAM_ERR;
    output [11:0] STAT_RX_DIAGWORD_INTFSTAT;
    output [11:0] STAT_RX_DIAGWORD_LANESTAT;
    output [255:0] STAT_RX_FC_STAT;
    output [11:0] STAT_RX_FRAMING_ERR;
    output STAT_RX_MEOP_ERR;
    output [11:0] STAT_RX_MF_ERR;
    output [11:0] STAT_RX_MF_LEN_ERR;
    output [11:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MSOP_ERR;
    output [7:0] STAT_RX_MUBITS;
    output STAT_RX_MUBITS_UPDATED;
    output STAT_RX_OVERFLOW_ERR;
    output STAT_RX_RETRANS_CRC24_ERR;
    output STAT_RX_RETRANS_DISC;
    output [15:0] STAT_RX_RETRANS_LATENCY;
    output STAT_RX_RETRANS_REQ;
    output STAT_RX_RETRANS_RETRY_ERR;
    output [7:0] STAT_RX_RETRANS_SEQ;
    output STAT_RX_RETRANS_SEQ_UPDATED;
    output [2:0] STAT_RX_RETRANS_STATE;
    output [4:0] STAT_RX_RETRANS_SUBSEQ;
    output STAT_RX_RETRANS_WDOG_ERR;
    output STAT_RX_RETRANS_WRAP_ERR;
    output [11:0] STAT_RX_SYNCED;
    output [11:0] STAT_RX_SYNCED_ERR;
    output [11:0] STAT_RX_WORD_SYNC;
    output STAT_TX_BURST_ERR;
    output STAT_TX_ERRINJ_BITERR_DONE;
    output STAT_TX_OVERFLOW_ERR;
    output STAT_TX_RETRANS_BURST_ERR;
    output STAT_TX_RETRANS_BUSY;
    output STAT_TX_RETRANS_RAM_PERROUT;
    output [8:0] STAT_TX_RETRANS_RAM_RADDR;
    output STAT_TX_RETRANS_RAM_RD_B0;
    output STAT_TX_RETRANS_RAM_RD_B1;
    output STAT_TX_RETRANS_RAM_RD_B2;
    output STAT_TX_RETRANS_RAM_RD_B3;
    output [1:0] STAT_TX_RETRANS_RAM_RSEL;
    output [8:0] STAT_TX_RETRANS_RAM_WADDR;
    output [643:0] STAT_TX_RETRANS_RAM_WDATA;
    output STAT_TX_RETRANS_RAM_WE_B0;
    output STAT_TX_RETRANS_RAM_WE_B1;
    output STAT_TX_RETRANS_RAM_WE_B2;
    output STAT_TX_RETRANS_RAM_WE_B3;
    output STAT_TX_UNDERFLOW_ERR;
    output TX_OVFOUT;
    output TX_RDYOUT;
    output [63:0] TX_SERDES_DATA00;
    output [63:0] TX_SERDES_DATA01;
    output [63:0] TX_SERDES_DATA02;
    output [63:0] TX_SERDES_DATA03;
    output [63:0] TX_SERDES_DATA04;
    output [63:0] TX_SERDES_DATA05;
    output [63:0] TX_SERDES_DATA06;
    output [63:0] TX_SERDES_DATA07;
    output [63:0] TX_SERDES_DATA08;
    output [63:0] TX_SERDES_DATA09;
    output [63:0] TX_SERDES_DATA10;
    output [63:0] TX_SERDES_DATA11;
    input CORE_CLK;
    input CTL_RX_FORCE_RESYNC;
    input CTL_RX_RETRANS_ACK;
    input CTL_RX_RETRANS_ENABLE;
    input CTL_RX_RETRANS_ERRIN;
    input CTL_RX_RETRANS_FORCE_REQ;
    input CTL_RX_RETRANS_RESET;
    input CTL_RX_RETRANS_RESET_MODE;
    input CTL_TX_DIAGWORD_INTFSTAT;
    input [11:0] CTL_TX_DIAGWORD_LANESTAT;
    input CTL_TX_ENABLE;
    input CTL_TX_ERRINJ_BITERR_GO;
    input [3:0] CTL_TX_ERRINJ_BITERR_LANE;
    input [255:0] CTL_TX_FC_STAT;
    input [7:0] CTL_TX_MUBITS;
    input CTL_TX_RETRANS_ENABLE;
    input CTL_TX_RETRANS_RAM_PERRIN;
    input [643:0] CTL_TX_RETRANS_RAM_RDATA;
    input CTL_TX_RETRANS_REQ;
    input CTL_TX_RETRANS_REQ_VALID;
    input [11:0] CTL_TX_RLIM_DELTA;
    input CTL_TX_RLIM_ENABLE;
    input [7:0] CTL_TX_RLIM_INTV;
    input [11:0] CTL_TX_RLIM_MAX;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input LBUS_CLK;
    input RX_BYPASS_FORCE_REALIGNIN;
    input RX_BYPASS_RDIN;
    input RX_RESET;
    input [11:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA00;
    input [63:0] RX_SERDES_DATA01;
    input [63:0] RX_SERDES_DATA02;
    input [63:0] RX_SERDES_DATA03;
    input [63:0] RX_SERDES_DATA04;
    input [63:0] RX_SERDES_DATA05;
    input [63:0] RX_SERDES_DATA06;
    input [63:0] RX_SERDES_DATA07;
    input [63:0] RX_SERDES_DATA08;
    input [63:0] RX_SERDES_DATA09;
    input [63:0] RX_SERDES_DATA10;
    input [63:0] RX_SERDES_DATA11;
    input [11:0] RX_SERDES_RESET;
    input TX_BCTLIN0;
    input TX_BCTLIN1;
    input TX_BCTLIN2;
    input TX_BCTLIN3;
    input [11:0] TX_BYPASS_CTRLIN;
    input [63:0] TX_BYPASS_DATAIN00;
    input [63:0] TX_BYPASS_DATAIN01;
    input [63:0] TX_BYPASS_DATAIN02;
    input [63:0] TX_BYPASS_DATAIN03;
    input [63:0] TX_BYPASS_DATAIN04;
    input [63:0] TX_BYPASS_DATAIN05;
    input [63:0] TX_BYPASS_DATAIN06;
    input [63:0] TX_BYPASS_DATAIN07;
    input [63:0] TX_BYPASS_DATAIN08;
    input [63:0] TX_BYPASS_DATAIN09;
    input [63:0] TX_BYPASS_DATAIN10;
    input [63:0] TX_BYPASS_DATAIN11;
    input TX_BYPASS_ENAIN;
    input [7:0] TX_BYPASS_GEARBOX_SEQIN;
    input [3:0] TX_BYPASS_MFRAMER_STATEIN;
    input [10:0] TX_CHANIN0;
    input [10:0] TX_CHANIN1;
    input [10:0] TX_CHANIN2;
    input [10:0] TX_CHANIN3;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input TX_RESET;
    input TX_SERDES_REFCLK;
    input TX_SERDES_REFCLK_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

