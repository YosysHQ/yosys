module a;
task to (
  input integer [3:0]x
);
endtask
endmodule

