module top();
endmodule
