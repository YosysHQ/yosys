module SLE (
	output Q,
	input ADn,
	input ALn,
	input CLK,
	input D,
	input LAT,
	input SD,
	input EN,
	input SLn
);
	reg q_latch, q_ff;

	always @(posedge CLK, negedge ALn) begin
		if (!ALn) begin
			q_ff <= !ADn;
		end else if (EN) begin
			if (!SLn)
				q_ff <= SD;
			else
				q_ff <= D;
		end
	end

	always @* begin
		if (!ALn) begin
			q_latch <= !ADn;
		end else if (CLK && EN) begin
			if (!SLn)
				q_ff <= SD;
			else
				q_ff <= D;
		end
	end

	assign Q = LAT ? q_latch : q_ff;
endmodule

module CFG1 (
	output O,
	input A
);
	parameter [1:0] INIT = 2'h0;
	assign O = INIT >> A;
endmodule

module CFG2 (
	output O,
	input A,
	input B
);
	parameter [3:0] INIT = 4'h0;
	assign O = INIT >> {B, A};
endmodule

module CFG3 (
	output O,
	input A,
	input B,
	input C
);
	parameter [7:0] INIT = 8'h0;
	assign O = INIT >> {C, B, A};
endmodule

module CFG4 (
	output O,
	input A,
	input B,
	input C,
	input D
);
	parameter [15:0] INIT = 16'h0;
	assign O = INIT >> {D, C, B, A};
endmodule
