/*
ISC License

Copyright (C) 2024 Microchip Technology Inc. and its subsidiaries

Permission to use, copy, modify, and/or distribute this software for any
purpose with or without fee is hereby granted, provided that the above
copyright notice and this permission notice appear in all copies.

THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
*/

module uram_sr(clk, wr, raddr, din, waddr, dout);
	input clk;
	input [11:0] din;
	input wr;
	input [5:0] waddr, raddr;
	output [11:0] dout;
	reg [5:0] raddr_reg;
	reg [11:0] mem [0:63];
	assign dout = mem[raddr_reg];

	integer i;
	initial begin
		for (i = 0; i < 64; i = i + 1) begin
			mem[i] = 12'hfff;
		end
	end

	always@(posedge clk) begin
		raddr_reg <= raddr; if(wr)
		mem[waddr]<= din;
	end
endmodule