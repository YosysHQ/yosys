module test(in, out);

input wire in;
output  out;
assign out = (in+in);
assign out = 74;
endmodule
