module x1_lev2(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, 
	pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, 
	pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, 
	pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, 
	pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, 
	pi50, po00, po01, po02, po03, po04, po05, po06, po07, po08, 
	po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, 
	po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, 
	po29, po30, po31, po32, po33, po34);

input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, 
	pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, 
	pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, 
	pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, 
	pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, 
	pi50;

output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, 
	po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, 
	po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, 
	po30, po31, po32, po33, po34;

wire po05, po16, po18, po24, po25, po28, po29, n270, n271, n272, 
	n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
	n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
	n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
	n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
	n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
	n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
	n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
	n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
	n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
	n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
	n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
	n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
	n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
	n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
	n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
	n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
	n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
	n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, 
	n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
	n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
	n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
	n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
	n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
	n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
	n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
	n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
	n533;

assign po05 = pi32;

assign po16 = pi37;

assign po18 = pi38;

assign po24 = pi23;

assign po25 = pi24;

assign po28 = pi48;

assign po29 = pi49;

  IV2 U294 ( .A(po32), .Z(po33));
  OR2 U295 ( .A(n270), .B(n271), .Z(po32));
  OR2 U296 ( .A(po25), .B(po05), .Z(n271));
  AN2 U297 ( .A(n272), .B(n273), .Z(n270));
  OR2 U298 ( .A(pi31), .B(po01), .Z(n273));
  AN2 U299 ( .A(n274), .B(pi18), .Z(po31));
  AN2 U300 ( .A(pi17), .B(n275), .Z(n274));
  AN2 U301 ( .A(n276), .B(n272), .Z(po30));
  OR2 U302 ( .A(n277), .B(n278), .Z(n276));
  AN2 U303 ( .A(n279), .B(n280), .Z(n278));
  OR2 U304 ( .A(n281), .B(pi31), .Z(n280));
  AN2 U305 ( .A(pi35), .B(n282), .Z(n281));
  AN2 U306 ( .A(n283), .B(n284), .Z(n277));
  OR2 U307 ( .A(n285), .B(n286), .Z(n284));
  AN2 U308 ( .A(pi31), .B(n287), .Z(n286));
  IV2 U309 ( .A(pi05), .Z(n287));
  AN2 U310 ( .A(n288), .B(pi35), .Z(n285));
  AN2 U311 ( .A(pi21), .B(pi13), .Z(n288));
  AN2 U312 ( .A(pi07), .B(n289), .Z(po27));
  OR2 U313 ( .A(n290), .B(n291), .Z(po26));
  OR2 U314 ( .A(n292), .B(n293), .Z(n291));
  AN2 U315 ( .A(n294), .B(n295), .Z(n293));
  AN2 U316 ( .A(n296), .B(n297), .Z(n295));
  AN2 U317 ( .A(pi33), .B(n298), .Z(n294));
  IV2 U318 ( .A(n299), .Z(n298));
  AN2 U319 ( .A(pi19), .B(pi00), .Z(n299));
  AN2 U320 ( .A(n300), .B(n301), .Z(n292));
  AN2 U321 ( .A(n302), .B(n303), .Z(n301));
  OR2 U322 ( .A(n304), .B(pi35), .Z(n303));
  AN2 U323 ( .A(n305), .B(pi25), .Z(n304));
  AN2 U324 ( .A(pi11), .B(n306), .Z(n305));
  AN2 U325 ( .A(n272), .B(n307), .Z(n302));
  AN2 U326 ( .A(n308), .B(pi01), .Z(n300));
  AN2 U327 ( .A(n279), .B(pi17), .Z(n308));
  AN2 U328 ( .A(pi34), .B(n309), .Z(n290));
  OR2 U329 ( .A(n310), .B(n311), .Z(po23));
  AN2 U330 ( .A(n312), .B(n313), .Z(n310));
  OR2 U331 ( .A(n314), .B(n315), .Z(po22));
  AN2 U332 ( .A(n316), .B(n317), .Z(n315));
  AN2 U333 ( .A(n318), .B(n319), .Z(n317));
  OR2 U334 ( .A(n320), .B(n272), .Z(n319));
  AN2 U335 ( .A(n321), .B(n322), .Z(n320));
  IV2 U336 ( .A(pi02), .Z(n322));
  AN2 U337 ( .A(n296), .B(n323), .Z(n321));
  OR2 U338 ( .A(pi09), .B(n324), .Z(n318));
  AN2 U339 ( .A(pi05), .B(pi21), .Z(n324));
  AN2 U340 ( .A(pi31), .B(n309), .Z(n316));
  AN2 U341 ( .A(n325), .B(n326), .Z(n314));
  AN2 U342 ( .A(n283), .B(n327), .Z(n325));
  OR2 U343 ( .A(n328), .B(n329), .Z(n327));
  OR2 U344 ( .A(n330), .B(n331), .Z(n329));
  OR2 U345 ( .A(n332), .B(n333), .Z(n331));
  AN2 U346 ( .A(po05), .B(n272), .Z(n333));
  AN2 U347 ( .A(pi43), .B(n296), .Z(n332));
  AN2 U348 ( .A(pi47), .B(pi39), .Z(n330));
  OR2 U349 ( .A(n334), .B(n335), .Z(n328));
  OR2 U350 ( .A(n336), .B(n337), .Z(n335));
  AN2 U351 ( .A(n338), .B(pi40), .Z(n337));
  AN2 U352 ( .A(n339), .B(n340), .Z(n338));
  AN2 U353 ( .A(n341), .B(n342), .Z(n336));
  AN2 U354 ( .A(n343), .B(n344), .Z(n342));
  AN2 U355 ( .A(n345), .B(pi41), .Z(n341));
  AN2 U356 ( .A(pi29), .B(n346), .Z(n334));
  OR2 U357 ( .A(n347), .B(n348), .Z(po21));
  AN2 U358 ( .A(pi09), .B(po05), .Z(n348));
  AN2 U359 ( .A(n349), .B(n350), .Z(n347));
  AN2 U360 ( .A(n346), .B(n279), .Z(n350));
  AN2 U361 ( .A(n351), .B(n326), .Z(n349));
  OR2 U362 ( .A(n352), .B(n353), .Z(po20));
  OR2 U363 ( .A(n354), .B(n355), .Z(n353));
  AN2 U364 ( .A(pi22), .B(po05), .Z(n355));
  AN2 U365 ( .A(n356), .B(n357), .Z(n354));
  OR2 U366 ( .A(n358), .B(n359), .Z(n356));
  OR2 U367 ( .A(po05), .B(n360), .Z(n359));
  AN2 U368 ( .A(n361), .B(n362), .Z(n360));
  OR2 U369 ( .A(n363), .B(n364), .Z(n362));
  AN2 U370 ( .A(n346), .B(n365), .Z(n364));
  AN2 U371 ( .A(n366), .B(pi14), .Z(n346));
  AN2 U372 ( .A(n367), .B(n343), .Z(n363));
  OR2 U373 ( .A(n368), .B(n365), .Z(n367));
  OR2 U374 ( .A(n351), .B(pi29), .Z(n365));
  AN2 U375 ( .A(pi28), .B(n345), .Z(n368));
  AN2 U376 ( .A(n309), .B(n369), .Z(n361));
  AN2 U377 ( .A(pi07), .B(n370), .Z(n358));
  OR2 U378 ( .A(pi28), .B(pi29), .Z(n370));
  OR2 U379 ( .A(n371), .B(n372), .Z(n352));
  AN2 U380 ( .A(pi01), .B(n373), .Z(n372));
  OR2 U381 ( .A(n374), .B(pi30), .Z(n373));
  AN2 U382 ( .A(pi10), .B(pi25), .Z(n374));
  AN2 U383 ( .A(n375), .B(n376), .Z(n371));
  OR2 U384 ( .A(pi40), .B(pi41), .Z(n376));
  OR2 U385 ( .A(n377), .B(n378), .Z(po19));
  OR2 U386 ( .A(n379), .B(n380), .Z(n378));
  AN2 U387 ( .A(pi42), .B(pi01), .Z(n380));
  AN2 U388 ( .A(pi12), .B(n381), .Z(n379));
  OR2 U389 ( .A(n382), .B(n383), .Z(n381));
  OR2 U390 ( .A(n384), .B(n385), .Z(n383));
  AN2 U391 ( .A(n386), .B(n369), .Z(n384));
  OR2 U392 ( .A(po34), .B(n387), .Z(n386));
  OR2 U393 ( .A(pi40), .B(pi26), .Z(n387));
  OR2 U394 ( .A(pi27), .B(pi28), .Z(po34));
  OR2 U395 ( .A(pi31), .B(pi29), .Z(n382));
  OR2 U396 ( .A(n388), .B(n389), .Z(n377));
  OR2 U397 ( .A(n390), .B(n391), .Z(n389));
  AN2 U398 ( .A(n392), .B(pi18), .Z(n391));
  AN2 U399 ( .A(pi17), .B(n393), .Z(n392));
  OR2 U400 ( .A(pi36), .B(pi40), .Z(n393));
  AN2 U401 ( .A(n394), .B(pi22), .Z(n390));
  AN2 U402 ( .A(n351), .B(n369), .Z(n394));
  AN2 U403 ( .A(pi00), .B(n395), .Z(n388));
  OR2 U404 ( .A(n396), .B(n397), .Z(n395));
  OR2 U405 ( .A(n385), .B(n398), .Z(n397));
  OR2 U406 ( .A(n399), .B(n400), .Z(n398));
  AN2 U407 ( .A(pi31), .B(n272), .Z(n399));
  OR2 U408 ( .A(n401), .B(n402), .Z(n385));
  OR2 U409 ( .A(pi41), .B(pi35), .Z(n402));
  OR2 U410 ( .A(po05), .B(pi43), .Z(n401));
  OR2 U411 ( .A(n403), .B(n404), .Z(n396));
  OR2 U412 ( .A(pi25), .B(n289), .Z(n404));
  OR2 U413 ( .A(pi34), .B(pi28), .Z(n403));
  IV2 U414 ( .A(po17), .Z(po15));
  OR2 U415 ( .A(n405), .B(n406), .Z(po17));
  OR2 U416 ( .A(n407), .B(n408), .Z(n406));
  OR2 U417 ( .A(n409), .B(n410), .Z(n408));
  AN2 U418 ( .A(pi28), .B(n411), .Z(n410));
  OR2 U419 ( .A(pi03), .B(n296), .Z(n411));
  AN2 U420 ( .A(n412), .B(n413), .Z(n409));
  OR2 U421 ( .A(n414), .B(n415), .Z(n413));
  AN2 U422 ( .A(pi02), .B(pi31), .Z(n415));
  AN2 U423 ( .A(n416), .B(n417), .Z(n414));
  AN2 U424 ( .A(n418), .B(n309), .Z(n416));
  OR2 U425 ( .A(pi25), .B(n272), .Z(n418));
  OR2 U426 ( .A(pi09), .B(n419), .Z(n412));
  AN2 U427 ( .A(n420), .B(n421), .Z(n419));
  AN2 U428 ( .A(n275), .B(n309), .Z(n421));
  OR2 U429 ( .A(pi25), .B(pi35), .Z(n275));
  AN2 U430 ( .A(n417), .B(pi21), .Z(n420));
  OR2 U431 ( .A(pi26), .B(n313), .Z(n407));
  AN2 U432 ( .A(pi33), .B(pi08), .Z(n313));
  OR2 U433 ( .A(n422), .B(n423), .Z(n405));
  OR2 U434 ( .A(po05), .B(pi27), .Z(n423));
  AN2 U435 ( .A(n424), .B(n425), .Z(po14));
  AN2 U436 ( .A(n426), .B(n309), .Z(n425));
  OR2 U437 ( .A(n427), .B(n428), .Z(n426));
  OR2 U438 ( .A(n429), .B(n430), .Z(n428));
  AN2 U439 ( .A(pi29), .B(n431), .Z(n430));
  OR2 U440 ( .A(pi43), .B(pi40), .Z(n427));
  AN2 U441 ( .A(n326), .B(pi07), .Z(n424));
  OR2 U442 ( .A(n432), .B(n433), .Z(po12));
  OR2 U443 ( .A(n434), .B(n435), .Z(n433));
  AN2 U444 ( .A(pi28), .B(n436), .Z(n435));
  OR2 U445 ( .A(n437), .B(pi21), .Z(n436));
  AN2 U446 ( .A(n438), .B(pi14), .Z(n437));
  AN2 U447 ( .A(n439), .B(n323), .Z(n438));
  OR2 U448 ( .A(n440), .B(n441), .Z(n439));
  IV2 U449 ( .A(n442), .Z(n441));
  AN2 U450 ( .A(n443), .B(pi15), .Z(n440));
  AN2 U451 ( .A(n444), .B(n445), .Z(n434));
  AN2 U452 ( .A(n446), .B(n312), .Z(n445));
  AN2 U453 ( .A(n447), .B(n448), .Z(n446));
  OR2 U454 ( .A(n282), .B(n307), .Z(n447));
  IV2 U455 ( .A(pi18), .Z(n307));
  AN2 U456 ( .A(n449), .B(pi40), .Z(n444));
  AN2 U457 ( .A(n450), .B(n451), .Z(n449));
  OR2 U458 ( .A(n339), .B(n297), .Z(n451));
  IV2 U459 ( .A(n452), .Z(n450));
  AN2 U460 ( .A(n453), .B(n339), .Z(n452));
  OR2 U461 ( .A(n340), .B(pi12), .Z(n453));
  AN2 U462 ( .A(pi02), .B(pi03), .Z(n340));
  AN2 U463 ( .A(pi46), .B(pi39), .Z(n432));
  IV2 U464 ( .A(po13), .Z(po11));
  OR2 U465 ( .A(n454), .B(n455), .Z(po13));
  OR2 U466 ( .A(n456), .B(n457), .Z(n455));
  AN2 U467 ( .A(pi25), .B(n458), .Z(n457));
  OR2 U468 ( .A(n459), .B(n460), .Z(n458));
  OR2 U469 ( .A(n461), .B(n462), .Z(n460));
  AN2 U470 ( .A(n463), .B(n464), .Z(n461));
  OR2 U471 ( .A(n282), .B(n465), .Z(n464));
  OR2 U472 ( .A(pi12), .B(pi09), .Z(n465));
  IV2 U473 ( .A(pi50), .Z(n463));
  AN2 U474 ( .A(pi07), .B(n466), .Z(n456));
  OR2 U475 ( .A(n467), .B(n468), .Z(n466));
  OR2 U476 ( .A(n469), .B(n429), .Z(n468));
  AN2 U477 ( .A(pi28), .B(n470), .Z(n429));
  AN2 U478 ( .A(n400), .B(n471), .Z(n469));
  OR2 U479 ( .A(pi40), .B(n431), .Z(n471));
  OR2 U480 ( .A(pi43), .B(n289), .Z(n467));
  AN2 U481 ( .A(pi19), .B(pi33), .Z(n289));
  OR2 U482 ( .A(po01), .B(n472), .Z(n454));
  OR2 U483 ( .A(po28), .B(po16), .Z(n472));
  OR2 U484 ( .A(n473), .B(n474), .Z(po10));
  AN2 U485 ( .A(n475), .B(pi41), .Z(n474));
  AN2 U486 ( .A(n476), .B(n477), .Z(n475));
  OR2 U487 ( .A(n297), .B(n343), .Z(n476));
  AN2 U488 ( .A(n478), .B(n479), .Z(n473));
  AN2 U489 ( .A(n283), .B(n296), .Z(n479));
  AN2 U490 ( .A(pi29), .B(n345), .Z(n478));
  IV2 U491 ( .A(n480), .Z(n345));
  IV2 U492 ( .A(po07), .Z(po09));
  OR2 U493 ( .A(n481), .B(n482), .Z(po08));
  AN2 U494 ( .A(pi45), .B(pi39), .Z(n482));
  AN2 U495 ( .A(n483), .B(n484), .Z(n481));
  OR2 U496 ( .A(n485), .B(n486), .Z(n484));
  AN2 U497 ( .A(pi29), .B(n312), .Z(n486));
  AN2 U498 ( .A(n296), .B(n309), .Z(n312));
  AN2 U499 ( .A(n351), .B(n487), .Z(n485));
  OR2 U500 ( .A(n488), .B(n326), .Z(n487));
  AN2 U501 ( .A(pi06), .B(n357), .Z(n488));
  AN2 U502 ( .A(pi03), .B(pi28), .Z(n351));
  AN2 U503 ( .A(n323), .B(n431), .Z(n483));
  OR2 U504 ( .A(n489), .B(n490), .Z(po07));
  OR2 U505 ( .A(pi33), .B(n311), .Z(n490));
  IV2 U506 ( .A(n491), .Z(n311));
  OR2 U507 ( .A(n492), .B(n493), .Z(n491));
  OR2 U508 ( .A(n494), .B(n297), .Z(n493));
  IV2 U509 ( .A(pi08), .Z(n297));
  AN2 U510 ( .A(n375), .B(n369), .Z(n494));
  IV2 U511 ( .A(n448), .Z(n375));
  OR2 U512 ( .A(n477), .B(n366), .Z(n448));
  OR2 U513 ( .A(n431), .B(n344), .Z(n477));
  IV2 U514 ( .A(pi16), .Z(n344));
  OR2 U515 ( .A(n495), .B(n496), .Z(n492));
  OR2 U516 ( .A(pi00), .B(n339), .Z(n496));
  AN2 U517 ( .A(n369), .B(n343), .Z(n339));
  IV2 U518 ( .A(n497), .Z(n495));
  OR2 U519 ( .A(n498), .B(pi40), .Z(n497));
  AN2 U520 ( .A(n369), .B(pi41), .Z(n498));
  OR2 U521 ( .A(po05), .B(n422), .Z(n489));
  OR2 U522 ( .A(po25), .B(po24), .Z(n422));
  OR2 U523 ( .A(n499), .B(n500), .Z(po06));
  AN2 U524 ( .A(pi27), .B(n501), .Z(n500));
  AN2 U525 ( .A(n502), .B(n503), .Z(n499));
  AN2 U526 ( .A(n504), .B(n480), .Z(n503));
  OR2 U527 ( .A(n431), .B(n366), .Z(n480));
  IV2 U528 ( .A(pi14), .Z(n431));
  AN2 U529 ( .A(n470), .B(n296), .Z(n504));
  IV2 U530 ( .A(pi07), .Z(n296));
  IV2 U531 ( .A(pi03), .Z(n470));
  AN2 U532 ( .A(pi28), .B(n279), .Z(n502));
  AN2 U533 ( .A(pi26), .B(n501), .Z(po04));
  OR2 U534 ( .A(pi21), .B(n323), .Z(n501));
  AN2 U535 ( .A(n505), .B(n506), .Z(po03));
  AN2 U536 ( .A(n507), .B(n279), .Z(n506));
  AN2 U537 ( .A(n369), .B(n283), .Z(n279));
  IV2 U538 ( .A(pi21), .Z(n369));
  AN2 U539 ( .A(n442), .B(n400), .Z(n507));
  OR2 U540 ( .A(pi29), .B(pi40), .Z(n400));
  OR2 U541 ( .A(n366), .B(n343), .Z(n442));
  IV2 U542 ( .A(pi06), .Z(n343));
  IV2 U543 ( .A(pi15), .Z(n366));
  AN2 U544 ( .A(n326), .B(pi14), .Z(n505));
  AN2 U545 ( .A(n508), .B(n443), .Z(n326));
  IV2 U546 ( .A(n357), .Z(n443));
  OR2 U547 ( .A(pi04), .B(pi20), .Z(n357));
  OR2 U548 ( .A(n509), .B(n510), .Z(po02));
  OR2 U549 ( .A(n511), .B(n512), .Z(n510));
  AN2 U550 ( .A(pi44), .B(pi39), .Z(n512));
  AN2 U551 ( .A(n513), .B(n514), .Z(n511));
  AN2 U552 ( .A(n515), .B(n516), .Z(n514));
  AN2 U553 ( .A(n309), .B(n306), .Z(n515));
  IV2 U554 ( .A(pi10), .Z(n306));
  AN2 U555 ( .A(n417), .B(pi25), .Z(n513));
  IV2 U556 ( .A(n517), .Z(n417));
  OR2 U557 ( .A(n518), .B(n519), .Z(n509));
  AN2 U558 ( .A(n520), .B(pi09), .Z(n519));
  AN2 U559 ( .A(n521), .B(pi02), .Z(n520));
  AN2 U560 ( .A(pi31), .B(n508), .Z(n521));
  IV2 U561 ( .A(pi22), .Z(n508));
  AN2 U562 ( .A(n522), .B(n272), .Z(n518));
  IV2 U563 ( .A(pi09), .Z(n272));
  AN2 U564 ( .A(n523), .B(n524), .Z(n522));
  AN2 U565 ( .A(n525), .B(pi35), .Z(n524));
  AN2 U566 ( .A(pi21), .B(n526), .Z(n525));
  IV2 U567 ( .A(pi13), .Z(n526));
  AN2 U568 ( .A(pi01), .B(n283), .Z(n523));
  AN2 U569 ( .A(n323), .B(n309), .Z(n283));
  IV2 U570 ( .A(pi00), .Z(n309));
  IV2 U571 ( .A(pi12), .Z(n323));
  OR2 U572 ( .A(n527), .B(n528), .Z(po00));
  AN2 U573 ( .A(po01), .B(n459), .Z(n528));
  OR2 U574 ( .A(pi30), .B(pi42), .Z(po01));
  AN2 U575 ( .A(pi25), .B(n529), .Z(n527));
  OR2 U576 ( .A(n530), .B(n517), .Z(n529));
  OR2 U577 ( .A(n531), .B(n532), .Z(n517));
  OR2 U578 ( .A(n462), .B(n459), .Z(n532));
  IV2 U579 ( .A(pi01), .Z(n459));
  IV2 U580 ( .A(pi11), .Z(n462));
  OR2 U581 ( .A(pi13), .B(pi12), .Z(n531));
  AN2 U582 ( .A(n533), .B(n282), .Z(n530));
  IV2 U583 ( .A(pi17), .Z(n282));
  IV2 U584 ( .A(n516), .Z(n533));
  OR2 U585 ( .A(pi09), .B(pi21), .Z(n516));

endmodule

module IV2(A,  Z);
  input A;
  output Z;

  assign Z = ~A;
endmodule

module AN2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A & B;
endmodule

module OR2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A | B;
endmodule
