module simple_assign (
    input wire in,
    output wire out
);

    assign out = in;

endmodule
