// ---------------------------------------

(* abc9_box_id=2 *)
module \$__ABC9_DPR16X4_COMB (input [3:0] A, S, output [3:0] Y);
endmodule
