module test;
endmodule
