module test(in, out);
input in;
output out;
parameter p = 10;

assign out = p;
endmodule
