module test(in, out, io);
inout io;
output out;
input in;

endmodule
