module TECH_AND18(input [17:0] in, output out);
assign out = &in;
endmodule

module TECH_AND4(input [3:0] in, output out);
assign out = &in;
endmodule
