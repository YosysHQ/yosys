module a(input wire x = 1'b0);
endmodule

