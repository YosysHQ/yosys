module C880_lev2(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, 
	pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, 
	pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, 
	pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, 
	pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, 
	pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, 
	po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, 
	po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, 
	po20, po21, po22, po23, po24, po25);

input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, 
	pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, 
	pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, 
	pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, 
	pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, 
	pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59;

output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, 
	po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, 
	po20, po21, po22, po23, po24, po25;

wire n137, n346, n364, n415, n295, n427, n351, n377, n454, n357, 
	n358, n359, n360, n361, n362, n363, n365, n366, n367, n368, 
	n369, n370, n371, n372, n373, n374, n375, n376, n378, n379, 
	n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
	n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
	n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
	n410, n411, n412, n413, n414, n416, n417, n418, n419, n420, 
	n421, n422, n423, n424, n425, n426, n428, n429, n430, n431, 
	n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
	n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
	n452, n453, n455, n456, n457, n458, n459, n460, n461, n462, 
	n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
	n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
	n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
	n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
	n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
	n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
	n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
	n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
	n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
	n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
	n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
	n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
	n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
	n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
	n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
	n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
	n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, 
	n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
	n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
	n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
	n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
	n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
	n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
	n693, n694, n695, n696;


assign po22 = n137;
assign po19 = n346;
assign po16 = n364;
assign po17 = n415;
assign po18 = n295;
assign po00 = n427;
assign po09 = n351;
assign po04 = n377;
assign po06 = n454;
  AN2 U371 ( .A(pi11), .B(pi08), .Z(n357));
  AN2 U372 ( .A(pi28), .B(n357), .Z(n346));
  AN2 U373 ( .A(pi41), .B(pi25), .Z(n369));
  AN2 U374 ( .A(pi52), .B(n369), .Z(n361));
  AN2 U375 ( .A(pi51), .B(pi54), .Z(n359));
  AN2 U376 ( .A(pi28), .B(pi31), .Z(n604));
  AN2 U377 ( .A(n604), .B(pi55), .Z(n358));
  AN2 U378 ( .A(n359), .B(n358), .Z(n602));
  AN2 U379 ( .A(pi53), .B(n602), .Z(n360));
  AN2 U380 ( .A(n361), .B(n360), .Z(n577));
  IV2 U381 ( .A(pi20), .Z(n607));
  OR2 U382 ( .A(n607), .B(pi25), .Z(n362));
  IV2 U383 ( .A(n362), .Z(n365));
  AN2 U384 ( .A(pi25), .B(n607), .Z(n363));
  OR2 U385 ( .A(n365), .B(n363), .Z(n367));
  AN2 U386 ( .A(pi41), .B(pi24), .Z(n378));
  AN2 U387 ( .A(n346), .B(n378), .Z(n366));
  AN2 U388 ( .A(n367), .B(n366), .Z(n373));
  AN2 U389 ( .A(pi28), .B(pi54), .Z(n368));
  AN2 U390 ( .A(pi20), .B(n368), .Z(n603));
  AN2 U391 ( .A(pi08), .B(n603), .Z(n371));
  IV2 U392 ( .A(pi56), .Z(n694));
  IV2 U393 ( .A(n369), .Z(n692));
  OR2 U394 ( .A(n694), .B(n692), .Z(n370));
  AN2 U395 ( .A(n371), .B(n370), .Z(n372));
  OR2 U396 ( .A(n373), .B(n372), .Z(n424));
  AN2 U397 ( .A(pi14), .B(n424), .Z(n384));
  AN2 U398 ( .A(pi56), .B(pi48), .Z(n608));
  AN2 U399 ( .A(n608), .B(n346), .Z(n374));
  AN2 U400 ( .A(pi07), .B(n374), .Z(n376));
  IV2 U401 ( .A(pi43), .Z(n375));
  AN2 U402 ( .A(n376), .B(n375), .Z(n406));
  AN2 U403 ( .A(pi20), .B(n406), .Z(n403));
  IV2 U404 ( .A(n378), .Z(n379));
  AN2 U405 ( .A(n346), .B(n379), .Z(n407));
  AN2 U406 ( .A(pi55), .B(n407), .Z(n399));
  AN2 U407 ( .A(pi44), .B(n399), .Z(n381));
  AN2 U408 ( .A(pi37), .B(pi54), .Z(n380));
  OR2 U409 ( .A(n381), .B(n380), .Z(n382));
  OR2 U410 ( .A(n403), .B(n382), .Z(n383));
  OR2 U411 ( .A(n384), .B(n383), .Z(n436));
  AN2 U412 ( .A(pi26), .B(n436), .Z(n385));
  OR2 U413 ( .A(n577), .B(n385), .Z(n386));
  AN2 U414 ( .A(pi34), .B(n386), .Z(n448));
  AN2 U415 ( .A(pi43), .B(pi05), .Z(n388));
  AN2 U416 ( .A(pi32), .B(n436), .Z(n387));
  OR2 U417 ( .A(n388), .B(n387), .Z(n446));
  AN2 U418 ( .A(pi08), .B(pi37), .Z(n393));
  AN2 U419 ( .A(pi50), .B(n399), .Z(n390));
  AN2 U420 ( .A(pi18), .B(n424), .Z(n389));
  OR2 U421 ( .A(n390), .B(n389), .Z(n391));
  OR2 U422 ( .A(n403), .B(n391), .Z(n392));
  OR2 U423 ( .A(n393), .B(n392), .Z(n494));
  AN2 U424 ( .A(pi27), .B(n494), .Z(n497));
  OR2 U425 ( .A(pi27), .B(n494), .Z(n499));
  AN2 U426 ( .A(pi20), .B(pi37), .Z(n398));
  AN2 U427 ( .A(pi45), .B(n399), .Z(n395));
  AN2 U428 ( .A(pi22), .B(n424), .Z(n394));
  OR2 U429 ( .A(n395), .B(n394), .Z(n396));
  OR2 U430 ( .A(n403), .B(n396), .Z(n397));
  OR2 U431 ( .A(n398), .B(n397), .Z(n536));
  AN2 U432 ( .A(pi17), .B(n536), .Z(n539));
  OR2 U433 ( .A(pi17), .B(n536), .Z(n541));
  AN2 U434 ( .A(pi23), .B(n424), .Z(n405));
  AN2 U435 ( .A(pi30), .B(pi37), .Z(n401));
  AN2 U436 ( .A(pi29), .B(n399), .Z(n400));
  OR2 U437 ( .A(n401), .B(n400), .Z(n402));
  OR2 U438 ( .A(n403), .B(n402), .Z(n404));
  OR2 U439 ( .A(n405), .B(n404), .Z(n579));
  AN2 U440 ( .A(pi21), .B(n579), .Z(n582));
  OR2 U441 ( .A(pi21), .B(n579), .Z(n584));
  AN2 U442 ( .A(n406), .B(pi55), .Z(n429));
  IV2 U443 ( .A(pi28), .Z(n409));
  AN2 U444 ( .A(n407), .B(pi20), .Z(n408));
  OR2 U445 ( .A(n409), .B(n408), .Z(n423));
  AN2 U446 ( .A(pi50), .B(n423), .Z(n411));
  AN2 U447 ( .A(pi42), .B(n424), .Z(n410));
  OR2 U448 ( .A(n411), .B(n410), .Z(n412));
  OR2 U449 ( .A(n429), .B(n412), .Z(n514));
  AN2 U450 ( .A(pi15), .B(n514), .Z(n517));
  OR2 U451 ( .A(pi15), .B(n514), .Z(n519));
  AN2 U452 ( .A(pi45), .B(n423), .Z(n414));
  AN2 U453 ( .A(pi40), .B(n424), .Z(n413));
  OR2 U454 ( .A(n414), .B(n413), .Z(n416));
  OR2 U455 ( .A(n429), .B(n416), .Z(n556));
  AN2 U456 ( .A(pi03), .B(n556), .Z(n559));
  OR2 U457 ( .A(pi03), .B(n556), .Z(n561));
  AN2 U458 ( .A(pi29), .B(n423), .Z(n418));
  AN2 U459 ( .A(pi04), .B(n424), .Z(n417));
  OR2 U460 ( .A(n418), .B(n417), .Z(n419));
  OR2 U461 ( .A(n429), .B(n419), .Z(n471));
  AN2 U462 ( .A(pi10), .B(n471), .Z(n480));
  OR2 U463 ( .A(pi10), .B(n471), .Z(n482));
  AN2 U464 ( .A(pi46), .B(n482), .Z(n420));
  OR2 U465 ( .A(n480), .B(n420), .Z(n562));
  AN2 U466 ( .A(n561), .B(n562), .Z(n421));
  OR2 U467 ( .A(n559), .B(n421), .Z(n520));
  AN2 U468 ( .A(n519), .B(n520), .Z(n422));
  OR2 U469 ( .A(n517), .B(n422), .Z(n449));
  AN2 U470 ( .A(pi44), .B(n423), .Z(n426));
  AN2 U471 ( .A(pi49), .B(n424), .Z(n425));
  OR2 U472 ( .A(n426), .B(n425), .Z(n428));
  OR2 U473 ( .A(n429), .B(n428), .Z(n464));
  AN2 U474 ( .A(n449), .B(n464), .Z(n432));
  OR2 U475 ( .A(n449), .B(n464), .Z(n430));
  AN2 U476 ( .A(pi09), .B(n430), .Z(n431));
  OR2 U477 ( .A(n432), .B(n431), .Z(n585));
  AN2 U478 ( .A(n584), .B(n585), .Z(n433));
  OR2 U479 ( .A(n582), .B(n433), .Z(n542));
  AN2 U480 ( .A(n541), .B(n542), .Z(n434));
  OR2 U481 ( .A(n539), .B(n434), .Z(n500));
  AN2 U482 ( .A(n499), .B(n500), .Z(n435));
  OR2 U483 ( .A(n497), .B(n435), .Z(n597));
  OR2 U484 ( .A(pi34), .B(n436), .Z(n598));
  AN2 U485 ( .A(n436), .B(pi34), .Z(n600));
  IV2 U486 ( .A(n600), .Z(n437));
  AN2 U487 ( .A(n598), .B(n437), .Z(n442));
  OR2 U488 ( .A(n597), .B(n442), .Z(n440));
  AN2 U489 ( .A(n597), .B(n442), .Z(n438));
  IV2 U490 ( .A(n438), .Z(n439));
  AN2 U491 ( .A(n440), .B(n439), .Z(n441));
  AN2 U492 ( .A(pi12), .B(n441), .Z(n444));
  AN2 U493 ( .A(n442), .B(pi19), .Z(n443));
  OR2 U494 ( .A(n444), .B(n443), .Z(n445));
  OR2 U495 ( .A(n446), .B(n445), .Z(n447));
  OR2 U496 ( .A(n448), .B(n447), .Z(n137));
  IV2 U497 ( .A(n464), .Z(n459));
  AN2 U498 ( .A(pi12), .B(n449), .Z(n456));
  AN2 U499 ( .A(n459), .B(n456), .Z(n453));
  IV2 U500 ( .A(n449), .Z(n450));
  AN2 U501 ( .A(n450), .B(pi12), .Z(n451));
  OR2 U502 ( .A(pi19), .B(n451), .Z(n458));
  AN2 U503 ( .A(n464), .B(n458), .Z(n452));
  OR2 U504 ( .A(n453), .B(n452), .Z(n455));
  IV2 U505 ( .A(pi09), .Z(n612));
  AN2 U506 ( .A(n455), .B(n612), .Z(n470));
  OR2 U507 ( .A(pi26), .B(n456), .Z(n457));
  AN2 U508 ( .A(n464), .B(n457), .Z(n462));
  AN2 U509 ( .A(n459), .B(n458), .Z(n460));
  OR2 U510 ( .A(n577), .B(n460), .Z(n461));
  OR2 U511 ( .A(n462), .B(n461), .Z(n463));
  AN2 U512 ( .A(pi09), .B(n463), .Z(n468));
  AN2 U513 ( .A(pi23), .B(pi05), .Z(n466));
  AN2 U514 ( .A(pi32), .B(n464), .Z(n465));
  OR2 U515 ( .A(n466), .B(n465), .Z(n467));
  OR2 U516 ( .A(n468), .B(n467), .Z(n469));
  OR2 U517 ( .A(n470), .B(n469), .Z(n295));
  AN2 U518 ( .A(pi26), .B(n480), .Z(n479));
  AN2 U519 ( .A(pi40), .B(pi05), .Z(n473));
  AN2 U520 ( .A(pi32), .B(n471), .Z(n472));
  OR2 U521 ( .A(n473), .B(n472), .Z(n477));
  AN2 U522 ( .A(pi38), .B(pi36), .Z(n475));
  AN2 U523 ( .A(pi10), .B(n577), .Z(n474));
  OR2 U524 ( .A(n475), .B(n474), .Z(n476));
  OR2 U525 ( .A(n477), .B(n476), .Z(n478));
  OR2 U526 ( .A(n479), .B(n478), .Z(n491));
  IV2 U527 ( .A(n480), .Z(n481));
  AN2 U528 ( .A(n482), .B(n481), .Z(n487));
  OR2 U529 ( .A(pi46), .B(n487), .Z(n485));
  AN2 U530 ( .A(pi46), .B(n487), .Z(n483));
  IV2 U531 ( .A(n483), .Z(n484));
  AN2 U532 ( .A(n485), .B(n484), .Z(n486));
  AN2 U533 ( .A(pi12), .B(n486), .Z(n489));
  AN2 U534 ( .A(n487), .B(pi19), .Z(n488));
  OR2 U535 ( .A(n489), .B(n488), .Z(n490));
  OR2 U536 ( .A(n491), .B(n490), .Z(n351));
  AN2 U537 ( .A(pi26), .B(n494), .Z(n492));
  OR2 U538 ( .A(n577), .B(n492), .Z(n493));
  AN2 U539 ( .A(pi27), .B(n493), .Z(n511));
  AN2 U540 ( .A(pi14), .B(pi05), .Z(n496));
  AN2 U541 ( .A(pi32), .B(n494), .Z(n495));
  OR2 U542 ( .A(n496), .B(n495), .Z(n509));
  IV2 U543 ( .A(n497), .Z(n498));
  AN2 U544 ( .A(n499), .B(n498), .Z(n505));
  OR2 U545 ( .A(n500), .B(n505), .Z(n503));
  AN2 U546 ( .A(n500), .B(n505), .Z(n501));
  IV2 U547 ( .A(n501), .Z(n502));
  AN2 U548 ( .A(n503), .B(n502), .Z(n504));
  AN2 U549 ( .A(pi12), .B(n504), .Z(n507));
  AN2 U550 ( .A(n505), .B(pi19), .Z(n506));
  OR2 U551 ( .A(n507), .B(n506), .Z(n508));
  OR2 U552 ( .A(n509), .B(n508), .Z(n510));
  OR2 U553 ( .A(n511), .B(n510), .Z(n364));
  AN2 U554 ( .A(pi26), .B(n514), .Z(n512));
  OR2 U555 ( .A(n577), .B(n512), .Z(n513));
  AN2 U556 ( .A(pi15), .B(n513), .Z(n533));
  AN2 U557 ( .A(pi49), .B(pi05), .Z(n531));
  AN2 U558 ( .A(pi33), .B(pi36), .Z(n516));
  AN2 U559 ( .A(pi32), .B(n514), .Z(n515));
  OR2 U560 ( .A(n516), .B(n515), .Z(n529));
  IV2 U561 ( .A(n517), .Z(n518));
  AN2 U562 ( .A(n519), .B(n518), .Z(n525));
  OR2 U563 ( .A(n520), .B(n525), .Z(n523));
  AN2 U564 ( .A(n520), .B(n525), .Z(n521));
  IV2 U565 ( .A(n521), .Z(n522));
  AN2 U566 ( .A(n523), .B(n522), .Z(n524));
  AN2 U567 ( .A(pi12), .B(n524), .Z(n527));
  AN2 U568 ( .A(n525), .B(pi19), .Z(n526));
  OR2 U569 ( .A(n527), .B(n526), .Z(n528));
  OR2 U570 ( .A(n529), .B(n528), .Z(n530));
  OR2 U571 ( .A(n531), .B(n530), .Z(n532));
  OR2 U572 ( .A(n533), .B(n532), .Z(n377));
  AN2 U573 ( .A(pi26), .B(n536), .Z(n534));
  OR2 U574 ( .A(n577), .B(n534), .Z(n535));
  AN2 U575 ( .A(pi17), .B(n535), .Z(n553));
  AN2 U576 ( .A(pi18), .B(pi05), .Z(n538));
  AN2 U577 ( .A(pi32), .B(n536), .Z(n537));
  OR2 U578 ( .A(n538), .B(n537), .Z(n551));
  IV2 U579 ( .A(n539), .Z(n540));
  AN2 U580 ( .A(n541), .B(n540), .Z(n547));
  OR2 U581 ( .A(n542), .B(n547), .Z(n545));
  AN2 U582 ( .A(n542), .B(n547), .Z(n543));
  IV2 U583 ( .A(n543), .Z(n544));
  AN2 U584 ( .A(n545), .B(n544), .Z(n546));
  AN2 U585 ( .A(pi12), .B(n546), .Z(n549));
  AN2 U586 ( .A(n547), .B(pi19), .Z(n548));
  OR2 U587 ( .A(n549), .B(n548), .Z(n550));
  OR2 U588 ( .A(n551), .B(n550), .Z(n552));
  OR2 U589 ( .A(n553), .B(n552), .Z(n415));
  AN2 U590 ( .A(pi26), .B(n556), .Z(n554));
  OR2 U591 ( .A(n577), .B(n554), .Z(n555));
  AN2 U592 ( .A(pi03), .B(n555), .Z(n575));
  AN2 U593 ( .A(pi42), .B(pi05), .Z(n573));
  AN2 U594 ( .A(pi47), .B(pi36), .Z(n558));
  AN2 U595 ( .A(pi32), .B(n556), .Z(n557));
  OR2 U596 ( .A(n558), .B(n557), .Z(n571));
  IV2 U597 ( .A(n559), .Z(n560));
  AN2 U598 ( .A(n561), .B(n560), .Z(n567));
  OR2 U599 ( .A(n562), .B(n567), .Z(n565));
  AN2 U600 ( .A(n562), .B(n567), .Z(n563));
  IV2 U601 ( .A(n563), .Z(n564));
  AN2 U602 ( .A(n565), .B(n564), .Z(n566));
  AN2 U603 ( .A(pi12), .B(n566), .Z(n569));
  AN2 U604 ( .A(n567), .B(pi19), .Z(n568));
  OR2 U605 ( .A(n569), .B(n568), .Z(n570));
  OR2 U606 ( .A(n571), .B(n570), .Z(n572));
  OR2 U607 ( .A(n573), .B(n572), .Z(n574));
  OR2 U608 ( .A(n575), .B(n574), .Z(n427));
  AN2 U609 ( .A(pi26), .B(n579), .Z(n576));
  OR2 U610 ( .A(n577), .B(n576), .Z(n578));
  AN2 U611 ( .A(pi21), .B(n578), .Z(n596));
  AN2 U612 ( .A(pi22), .B(pi05), .Z(n581));
  AN2 U613 ( .A(pi32), .B(n579), .Z(n580));
  OR2 U614 ( .A(n581), .B(n580), .Z(n594));
  IV2 U615 ( .A(n582), .Z(n583));
  AN2 U616 ( .A(n584), .B(n583), .Z(n590));
  OR2 U617 ( .A(n585), .B(n590), .Z(n588));
  AN2 U618 ( .A(n585), .B(n590), .Z(n586));
  IV2 U619 ( .A(n586), .Z(n587));
  AN2 U620 ( .A(n588), .B(n587), .Z(n589));
  AN2 U621 ( .A(pi12), .B(n589), .Z(n592));
  AN2 U622 ( .A(n590), .B(pi19), .Z(n591));
  OR2 U623 ( .A(n592), .B(n591), .Z(n593));
  OR2 U624 ( .A(n594), .B(n593), .Z(n595));
  OR2 U625 ( .A(n596), .B(n595), .Z(n454));
  AN2 U626 ( .A(n598), .B(n597), .Z(n599));
  OR2 U627 ( .A(n600), .B(n599), .Z(po07));
  OR2 U628 ( .A(pi58), .B(pi00), .Z(n609));
  AN2 U629 ( .A(pi59), .B(n609), .Z(po24));
  AN2 U630 ( .A(n602), .B(pi57), .Z(n601));
  AN2 U631 ( .A(pi41), .B(n601), .Z(po13));
  AN2 U632 ( .A(pi48), .B(n602), .Z(po08));
  AN2 U633 ( .A(n603), .B(pi31), .Z(po03));
  AN2 U634 ( .A(pi48), .B(pi16), .Z(n610));
  AN2 U635 ( .A(pi25), .B(n610), .Z(po25));
  AN2 U636 ( .A(pi11), .B(n604), .Z(n605));
  IV2 U637 ( .A(n605), .Z(n606));
  OR2 U638 ( .A(n607), .B(n606), .Z(n691));
  OR2 U639 ( .A(po25), .B(n691), .Z(po02));
  AN2 U640 ( .A(n608), .B(pi25), .Z(po10));
  AN2 U641 ( .A(pi13), .B(n609), .Z(po12));
  AN2 U642 ( .A(pi07), .B(n610), .Z(po14));
  IV2 U643 ( .A(pi15), .Z(n611));
  AN2 U644 ( .A(pi09), .B(n611), .Z(n614));
  AN2 U645 ( .A(pi15), .B(n612), .Z(n613));
  OR2 U646 ( .A(n614), .B(n613), .Z(n618));
  IV2 U647 ( .A(pi35), .Z(n654));
  OR2 U648 ( .A(n654), .B(pi06), .Z(n617));
  IV2 U649 ( .A(pi06), .Z(n615));
  OR2 U650 ( .A(n615), .B(pi35), .Z(n616));
  AN2 U651 ( .A(n617), .B(n616), .Z(n619));
  OR2 U652 ( .A(n618), .B(n619), .Z(n622));
  AN2 U653 ( .A(n619), .B(n618), .Z(n620));
  IV2 U654 ( .A(n620), .Z(n621));
  AN2 U655 ( .A(n622), .B(n621), .Z(n628));
  IV2 U656 ( .A(pi10), .Z(n624));
  OR2 U657 ( .A(n624), .B(pi03), .Z(n623));
  IV2 U658 ( .A(n623), .Z(n626));
  AN2 U659 ( .A(pi03), .B(n624), .Z(n625));
  OR2 U660 ( .A(n626), .B(n625), .Z(n627));
  OR2 U661 ( .A(n628), .B(n627), .Z(n631));
  AN2 U662 ( .A(n628), .B(n627), .Z(n629));
  IV2 U663 ( .A(n629), .Z(n630));
  AN2 U664 ( .A(n631), .B(n630), .Z(n637));
  IV2 U665 ( .A(pi34), .Z(n632));
  AN2 U666 ( .A(pi27), .B(n632), .Z(n635));
  OR2 U667 ( .A(n632), .B(pi27), .Z(n633));
  IV2 U668 ( .A(n633), .Z(n634));
  OR2 U669 ( .A(n635), .B(n634), .Z(n636));
  OR2 U670 ( .A(n637), .B(n636), .Z(n640));
  AN2 U671 ( .A(n637), .B(n636), .Z(n638));
  IV2 U672 ( .A(n638), .Z(n639));
  AN2 U673 ( .A(n640), .B(n639), .Z(n647));
  IV2 U674 ( .A(pi21), .Z(n642));
  OR2 U675 ( .A(n642), .B(pi17), .Z(n641));
  IV2 U676 ( .A(n641), .Z(n644));
  AN2 U677 ( .A(pi17), .B(n642), .Z(n643));
  OR2 U678 ( .A(n644), .B(n643), .Z(n646));
  OR2 U679 ( .A(n647), .B(n646), .Z(n645));
  IV2 U680 ( .A(n645), .Z(n649));
  AN2 U681 ( .A(n647), .B(n646), .Z(n648));
  OR2 U682 ( .A(n649), .B(n648), .Z(po15));
  IV2 U683 ( .A(pi42), .Z(n650));
  AN2 U684 ( .A(pi49), .B(n650), .Z(n653));
  IV2 U685 ( .A(pi49), .Z(n651));
  AN2 U686 ( .A(pi42), .B(n651), .Z(n652));
  OR2 U687 ( .A(n653), .B(n652), .Z(n658));
  OR2 U688 ( .A(n654), .B(pi39), .Z(n657));
  IV2 U689 ( .A(pi39), .Z(n655));
  OR2 U690 ( .A(n655), .B(pi35), .Z(n656));
  AN2 U691 ( .A(n657), .B(n656), .Z(n659));
  OR2 U692 ( .A(n658), .B(n659), .Z(n662));
  AN2 U693 ( .A(n659), .B(n658), .Z(n660));
  IV2 U694 ( .A(n660), .Z(n661));
  AN2 U695 ( .A(n662), .B(n661), .Z(n668));
  IV2 U696 ( .A(pi04), .Z(n664));
  OR2 U697 ( .A(n664), .B(pi18), .Z(n663));
  IV2 U698 ( .A(n663), .Z(n666));
  AN2 U699 ( .A(pi18), .B(n664), .Z(n665));
  OR2 U700 ( .A(n666), .B(n665), .Z(n667));
  OR2 U701 ( .A(n668), .B(n667), .Z(n671));
  AN2 U702 ( .A(n668), .B(n667), .Z(n669));
  IV2 U703 ( .A(n669), .Z(n670));
  AN2 U704 ( .A(n671), .B(n670), .Z(n677));
  IV2 U705 ( .A(pi22), .Z(n673));
  OR2 U706 ( .A(n673), .B(pi14), .Z(n672));
  IV2 U707 ( .A(n672), .Z(n675));
  AN2 U708 ( .A(pi14), .B(n673), .Z(n674));
  OR2 U709 ( .A(n675), .B(n674), .Z(n676));
  OR2 U710 ( .A(n677), .B(n676), .Z(n680));
  AN2 U711 ( .A(n677), .B(n676), .Z(n678));
  IV2 U712 ( .A(n678), .Z(n679));
  AN2 U713 ( .A(n680), .B(n679), .Z(n687));
  IV2 U714 ( .A(pi40), .Z(n682));
  OR2 U715 ( .A(n682), .B(pi23), .Z(n681));
  IV2 U716 ( .A(n681), .Z(n684));
  AN2 U717 ( .A(pi23), .B(n682), .Z(n683));
  OR2 U718 ( .A(n684), .B(n683), .Z(n686));
  OR2 U719 ( .A(n687), .B(n686), .Z(n685));
  IV2 U720 ( .A(n685), .Z(n689));
  AN2 U721 ( .A(n687), .B(n686), .Z(n688));
  OR2 U722 ( .A(n689), .B(n688), .Z(po20));
  AN2 U723 ( .A(pi01), .B(pi02), .Z(po21));
  IV2 U724 ( .A(po25), .Z(n690));
  OR2 U725 ( .A(n691), .B(n690), .Z(po23));
  IV2 U726 ( .A(pi16), .Z(n696));
  OR2 U727 ( .A(n692), .B(n696), .Z(po11));
  AN2 U728 ( .A(pi07), .B(pi41), .Z(n693));
  IV2 U729 ( .A(n693), .Z(n695));
  OR2 U730 ( .A(n694), .B(n695), .Z(po01));
  OR2 U731 ( .A(n696), .B(n695), .Z(po05));

endmodule

module IV2(A,  Z);
  input A;
  output Z;

  assign Z = ~A;
endmodule

module AN2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A & B;
endmodule

module OR2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A | B;
endmodule
