module TECH_OR18(input [17:0] in, output out);
assign out = |in;
endmodule

module TECH_OR4(input [3:0] in, output out);
assign out = |in;
endmodule
