module test(in1, in2, out1, out2, io1, io2);
inout [1:0] io1;
inout [0:1] io2;
output [1:0] out1;
output [0:1] out2;
input [1:0] in1;
input [0:1] in2;

endmodule
