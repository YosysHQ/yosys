module a;
task to (
  input [3]x
);
endtask
endmodule

