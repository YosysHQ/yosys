module undriven_replay (
	input wire in,
	output wire out,
	output wire undrv
);
	assign out = in;
endmodule
