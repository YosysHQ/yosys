module test(output out, input in);

assign out = +in;
endmodule
