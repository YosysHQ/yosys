module sv_top(input logic a, output logic y);
	assign y = a;
endmodule
