(* blackbox *)
module NX_BD(I, O);
    input I;
    output O;
    parameter mode = "global_lowskew";
endmodule

(* blackbox *)
module NX_BFF(I, O);
    input I;
    output O;
endmodule

(* blackbox *)
module NX_BFR(I, O);
    input I;
    output O;
    parameter data_inv = 1'b0;
    parameter iobname = "";
    parameter location = "";
    parameter mode = 0;
    parameter path = 0;
    parameter ring = 0;
endmodule

//(* blackbox *)
//module NX_CY(A1, A2, A3, A4, B1, B2, B3, B4, CI, CO, S1, S2, S3, S4);
//    input A1;
//    input A2;
//    input A3;
//    input A4;
//    input B1;
//    input B2;
//    input B3;
//    input B4;
//    input CI;
//    output CO;
//    output S1;
//    output S2;
//    output S3;
//    output S4;
//    parameter add_carry = 0;
//endmodule

(* blackbox *)
module NX_DES(FCK, SCK, R, IO, DCK, DRL, DIG, FZ, FLD, FLG, O, DS, DRA, DRI, DRO, DID);
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    input FCK;
    output FLD;
    output FLG;
    input FZ;
    input IO;
    output [4:0] O;
    input R;
    input SCK;
    parameter data_size = 5;
    parameter differential = "";
    parameter dpath_dynamic = 1'b0;
    parameter drive = "";
    parameter inputDelayLine = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

//(* blackbox *)
//module NX_DFF(I, CK, L, R, O);
//    input CK;
//    input I;
//    input L;
//    output O;
//    input R;
//    parameter dff_ctxt = 1'b0;
//    parameter dff_edge = 1'b0;
//    parameter dff_init = 1'b0;
//    parameter dff_load = 1'b0;
//    parameter dff_sync = 1'b0;
//    parameter dff_type = 1'b0;
//endmodule

(* blackbox *)
module NX_DFR(I, CK, L, R, O);
    input CK;
    input I;
    input L;
    output O;
    input R;
    parameter data_inv = 1'b0;
    parameter dff_edge = 1'b0;
    parameter dff_init = 1'b0;
    parameter dff_load = 1'b0;
    parameter dff_sync = 1'b0;
    parameter dff_type = 1'b0;
    parameter iobname = "";
    parameter location = "";
    parameter mode = 0;
    parameter path = 0;
    parameter ring = 0;
endmodule

(* blackbox *)
module NX_ECC(CKD, CHK, COR, ERR);
    input CHK;
    input CKD;
    output COR;
    output ERR;
endmodule

(* blackbox *)
module NX_HSSL_L_FULL(hssl_clk_user_i, hssl_clk_ref_i, hssl_clock_o, usr_com_tx_pma_pre_sign_i, usr_com_tx_pma_pre_en_i, usr_com_tx_pma_main_sign_i, usr_com_rx_pma_m_eye_i, usr_com_tx_pma_post_sign_i, usr_pll_pma_rst_n_i, usr_main_rst_n_i, usr_calibrate_pma_en_i, usr_pcs_ctrl_pll_lock_en_i, usr_pcs_ctrl_ovs_en_i, usr_pll_lock_o, usr_calibrate_pma_out_o, pma_clk_ext_i, usr_tx0_ctrl_replace_en_i, usr_tx0_rst_n_i, usr_tx0_pma_clk_en_i, usr_tx0_busy_o, pma_tx0_o
, usr_rx0_ctrl_dscr_en_i, usr_rx0_ctrl_dec_en_i, usr_rx0_ctrl_align_en_i, usr_rx0_ctrl_align_sync_i, usr_rx0_ctrl_replace_en_i, usr_rx0_ctrl_el_buff_rst_i, usr_rx0_ctrl_el_buff_fifo_en_i, usr_rx0_rst_n_i, usr_rx0_pma_cdr_rst_i, usr_rx0_pma_ckgen_rst_n_i, usr_rx0_pma_pll_rst_n_i, usr_rx0_pma_loss_of_signal_o, usr_rx0_ctrl_char_is_aligned_o, usr_rx0_busy_o, usr_rx0_pll_lock_o, pma_rx0_i, usr_tx1_ctrl_replace_en_i, usr_tx1_rst_n_i, usr_tx1_pma_clk_en_i, usr_tx1_busy_o, pma_tx1_o
, usr_rx1_ctrl_dscr_en_i, usr_rx1_ctrl_dec_en_i, usr_rx1_ctrl_align_en_i, usr_rx1_ctrl_align_sync_i, usr_rx1_ctrl_replace_en_i, usr_rx1_ctrl_el_buff_rst_i, usr_rx1_ctrl_el_buff_fifo_en_i, usr_rx1_rst_n_i, usr_rx1_pma_cdr_rst_i, usr_rx1_pma_ckgen_rst_n_i, usr_rx1_pma_pll_rst_n_i, usr_rx1_pma_loss_of_signal_o, usr_rx1_ctrl_char_is_aligned_o, usr_rx1_busy_o, usr_rx1_pll_lock_o, pma_rx1_i, usr_tx2_ctrl_replace_en_i, usr_tx2_rst_n_i, usr_tx2_pma_clk_en_i, usr_tx2_busy_o, pma_tx2_o
, usr_rx2_ctrl_dscr_en_i, usr_rx2_ctrl_dec_en_i, usr_rx2_ctrl_align_en_i, usr_rx2_ctrl_align_sync_i, usr_rx2_ctrl_replace_en_i, usr_rx2_ctrl_el_buff_rst_i, usr_rx2_ctrl_el_buff_fifo_en_i, usr_rx2_rst_n_i, usr_rx2_pma_cdr_rst_i, usr_rx2_pma_ckgen_rst_n_i, usr_rx2_pma_pll_rst_n_i, usr_rx2_pma_loss_of_signal_o, usr_rx2_ctrl_char_is_aligned_o, usr_rx2_busy_o, usr_rx2_pll_lock_o, pma_rx2_i, usr_tx3_ctrl_replace_en_i, usr_tx3_rst_n_i, usr_tx3_pma_clk_en_i, usr_tx3_busy_o, pma_tx3_o
, usr_rx3_ctrl_dscr_en_i, usr_rx3_ctrl_dec_en_i, usr_rx3_ctrl_align_en_i, usr_rx3_ctrl_align_sync_i, usr_rx3_ctrl_replace_en_i, usr_rx3_ctrl_el_buff_rst_i, usr_rx3_ctrl_el_buff_fifo_en_i, usr_rx3_rst_n_i, usr_rx3_pma_cdr_rst_i, usr_rx3_pma_ckgen_rst_n_i, usr_rx3_pma_pll_rst_n_i, usr_rx3_pma_loss_of_signal_o, usr_rx3_ctrl_char_is_aligned_o, usr_rx3_busy_o, usr_rx3_pll_lock_o, pma_rx3_i, usr_tx4_ctrl_replace_en_i, usr_tx4_rst_n_i, usr_tx4_pma_clk_en_i, usr_tx4_busy_o, pma_tx4_o
, usr_rx4_ctrl_dscr_en_i, usr_rx4_ctrl_dec_en_i, usr_rx4_ctrl_align_en_i, usr_rx4_ctrl_align_sync_i, usr_rx4_ctrl_replace_en_i, usr_rx4_ctrl_el_buff_rst_i, usr_rx4_ctrl_el_buff_fifo_en_i, usr_rx4_rst_n_i, usr_rx4_pma_cdr_rst_i, usr_rx4_pma_ckgen_rst_n_i, usr_rx4_pma_pll_rst_n_i, usr_rx4_pma_loss_of_signal_o, usr_rx4_ctrl_char_is_aligned_o, usr_rx4_busy_o, usr_rx4_pll_lock_o, pma_rx4_i, usr_tx5_ctrl_replace_en_i, usr_tx5_rst_n_i, usr_tx5_pma_clk_en_i, usr_tx5_busy_o, pma_tx5_o
, usr_rx5_ctrl_dscr_en_i, usr_rx5_ctrl_dec_en_i, usr_rx5_ctrl_align_en_i, usr_rx5_ctrl_align_sync_i, usr_rx5_ctrl_replace_en_i, usr_rx5_ctrl_el_buff_rst_i, usr_rx5_ctrl_el_buff_fifo_en_i, usr_rx5_rst_n_i, usr_rx5_pma_cdr_rst_i, usr_rx5_pma_ckgen_rst_n_i, usr_rx5_pma_pll_rst_n_i, usr_rx5_pma_loss_of_signal_o, usr_rx5_ctrl_char_is_aligned_o, usr_rx5_busy_o, usr_rx5_pll_lock_o, pma_rx5_i, usr_com_tx_pma_main_en_i, usr_com_tx_pma_margin_sel_i, usr_com_tx_pma_margin_input_sel_i, usr_com_tx_pma_margin_sel_var_i, usr_com_tx_pma_margin_input_sel_var_i
, usr_com_tx_pma_post_en_i, usr_com_tx_pma_post_input_sel_i, usr_com_tx_pma_post_input_sel_var_i, usr_com_rx_pma_ctle_cap_i, usr_com_rx_pma_ctle_resp_i, usr_com_rx_pma_ctle_resn_i, usr_com_ctrl_tx_sel_i, usr_com_ctrl_rx_sel_i, usr_calibrate_pma_res_p1_i, usr_calibrate_pma_res_n2_i, usr_calibrate_pma_res_n3_i, usr_calibrate_pma_res_p4_i, usr_calibrate_pma_sel_i, usr_main_test_i, usr_main_test_o, usr_tx0_ctrl_enc_en_i, usr_tx0_ctrl_char_is_k_i, usr_tx0_ctrl_scr_en_i, usr_tx0_ctrl_end_of_multiframe_i, usr_tx0_ctrl_end_of_frame_i, usr_tx0_test_i
, usr_tx0_data_i, usr_tx0_test_o, usr_rx0_data_o, usr_rx0_ctrl_ovs_bit_sel_i, usr_rx0_test_i, usr_rx0_ctrl_char_is_comma_o, usr_rx0_ctrl_char_is_k_o, usr_rx0_ctrl_not_in_table_o, usr_rx0_ctrl_disp_err_o, usr_rx0_ctrl_char_is_a_o, usr_rx0_ctrl_char_is_f_o, usr_rx0_test_o, usr_tx1_ctrl_enc_en_i, usr_tx1_ctrl_char_is_k_i, usr_tx1_ctrl_scr_en_i, usr_tx1_ctrl_end_of_multiframe_i, usr_tx1_ctrl_end_of_frame_i, usr_tx1_test_i, usr_tx1_data_i, usr_tx1_test_o, usr_rx1_data_o
, usr_rx1_ctrl_ovs_bit_sel_i, usr_rx1_test_i, usr_rx1_ctrl_char_is_comma_o, usr_rx1_ctrl_char_is_k_o, usr_rx1_ctrl_not_in_table_o, usr_rx1_ctrl_disp_err_o, usr_rx1_ctrl_char_is_a_o, usr_rx1_ctrl_char_is_f_o, usr_rx1_test_o, usr_tx2_ctrl_enc_en_i, usr_tx2_ctrl_char_is_k_i, usr_tx2_ctrl_scr_en_i, usr_tx2_ctrl_end_of_multiframe_i, usr_tx2_ctrl_end_of_frame_i, usr_tx2_test_i, usr_tx2_data_i, usr_tx2_test_o, usr_rx2_data_o, usr_rx2_ctrl_ovs_bit_sel_i, usr_rx2_test_i, usr_rx2_ctrl_char_is_comma_o
, usr_rx2_ctrl_char_is_k_o, usr_rx2_ctrl_not_in_table_o, usr_rx2_ctrl_disp_err_o, usr_rx2_ctrl_char_is_a_o, usr_rx2_ctrl_char_is_f_o, usr_rx2_test_o, usr_tx3_ctrl_enc_en_i, usr_tx3_ctrl_char_is_k_i, usr_tx3_ctrl_scr_en_i, usr_tx3_ctrl_end_of_multiframe_i, usr_tx3_ctrl_end_of_frame_i, usr_tx3_test_i, usr_tx3_data_i, usr_tx3_test_o, usr_rx3_data_o, usr_rx3_ctrl_ovs_bit_sel_i, usr_rx3_test_i, usr_rx3_ctrl_char_is_comma_o, usr_rx3_ctrl_char_is_k_o, usr_rx3_ctrl_not_in_table_o, usr_rx3_ctrl_disp_err_o
, usr_rx3_ctrl_char_is_a_o, usr_rx3_ctrl_char_is_f_o, usr_rx3_test_o, usr_tx4_ctrl_enc_en_i, usr_tx4_ctrl_char_is_k_i, usr_tx4_ctrl_scr_en_i, usr_tx4_ctrl_end_of_multiframe_i, usr_tx4_ctrl_end_of_frame_i, usr_tx4_test_i, usr_tx4_data_i, usr_tx4_test_o, usr_rx4_data_o, usr_rx4_ctrl_ovs_bit_sel_i, usr_rx4_test_i, usr_rx4_ctrl_char_is_comma_o, usr_rx4_ctrl_char_is_k_o, usr_rx4_ctrl_not_in_table_o, usr_rx4_ctrl_disp_err_o, usr_rx4_ctrl_char_is_a_o, usr_rx4_ctrl_char_is_f_o, usr_rx4_test_o
, usr_tx5_ctrl_enc_en_i, usr_tx5_ctrl_char_is_k_i, usr_tx5_ctrl_scr_en_i, usr_tx5_ctrl_end_of_multiframe_i, usr_tx5_ctrl_end_of_frame_i, usr_tx5_test_i, usr_tx5_data_i, usr_tx5_test_o, usr_rx5_data_o, usr_rx5_ctrl_ovs_bit_sel_i, usr_rx5_test_i, usr_rx5_ctrl_char_is_comma_o, usr_rx5_ctrl_char_is_k_o, usr_rx5_ctrl_not_in_table_o, usr_rx5_ctrl_disp_err_o, usr_rx5_ctrl_char_is_a_o, usr_rx5_ctrl_char_is_f_o, usr_rx5_test_o, usr_com_tx_pma_pre_input_sel_i);
    input hssl_clk_ref_i;
    input hssl_clk_user_i;
    output hssl_clock_o;
    input pma_clk_ext_i;
    input pma_rx0_i;
    input pma_rx1_i;
    input pma_rx2_i;
    input pma_rx3_i;
    input pma_rx4_i;
    input pma_rx5_i;
    output pma_tx0_o;
    output pma_tx1_o;
    output pma_tx2_o;
    output pma_tx3_o;
    output pma_tx4_o;
    output pma_tx5_o;
    input usr_calibrate_pma_en_i;
    output usr_calibrate_pma_out_o;
    input [7:0] usr_calibrate_pma_res_n2_i;
    input [7:0] usr_calibrate_pma_res_n3_i;
    input [7:0] usr_calibrate_pma_res_p1_i;
    input [7:0] usr_calibrate_pma_res_p4_i;
    input [3:0] usr_calibrate_pma_sel_i;
    input [5:0] usr_com_ctrl_rx_sel_i;
    input [5:0] usr_com_ctrl_tx_sel_i;
    input [3:0] usr_com_rx_pma_ctle_cap_i;
    input [3:0] usr_com_rx_pma_ctle_resn_i;
    input [3:0] usr_com_rx_pma_ctle_resp_i;
    input usr_com_rx_pma_m_eye_i;
    input [5:0] usr_com_tx_pma_main_en_i;
    input usr_com_tx_pma_main_sign_i;
    input [3:0] usr_com_tx_pma_margin_input_sel_i;
    input [4:0] usr_com_tx_pma_margin_input_sel_var_i;
    input [3:0] usr_com_tx_pma_margin_sel_i;
    input [4:0] usr_com_tx_pma_margin_sel_var_i;
    input [4:0] usr_com_tx_pma_post_en_i;
    input [3:0] usr_com_tx_pma_post_input_sel_i;
    input [3:0] usr_com_tx_pma_post_input_sel_var_i;
    input usr_com_tx_pma_post_sign_i;
    input usr_com_tx_pma_pre_en_i;
    input [3:0] usr_com_tx_pma_pre_input_sel_i;
    input usr_com_tx_pma_pre_sign_i;
    input usr_main_rst_n_i;
    input [7:0] usr_main_test_i;
    output [7:0] usr_main_test_o;
    input usr_pcs_ctrl_ovs_en_i;
    input usr_pcs_ctrl_pll_lock_en_i;
    output usr_pll_lock_o;
    input usr_pll_pma_rst_n_i;
    output usr_rx0_busy_o;
    input usr_rx0_ctrl_align_en_i;
    input usr_rx0_ctrl_align_sync_i;
    output [7:0] usr_rx0_ctrl_char_is_a_o;
    output usr_rx0_ctrl_char_is_aligned_o;
    output [7:0] usr_rx0_ctrl_char_is_comma_o;
    output [7:0] usr_rx0_ctrl_char_is_f_o;
    output [7:0] usr_rx0_ctrl_char_is_k_o;
    input usr_rx0_ctrl_dec_en_i;
    output [7:0] usr_rx0_ctrl_disp_err_o;
    input usr_rx0_ctrl_dscr_en_i;
    input usr_rx0_ctrl_el_buff_fifo_en_i;
    input usr_rx0_ctrl_el_buff_rst_i;
    output [7:0] usr_rx0_ctrl_not_in_table_o;
    input [1:0] usr_rx0_ctrl_ovs_bit_sel_i;
    input usr_rx0_ctrl_replace_en_i;
    output [63:0] usr_rx0_data_o;
    output usr_rx0_pll_lock_o;
    input usr_rx0_pma_cdr_rst_i;
    input usr_rx0_pma_ckgen_rst_n_i;
    output usr_rx0_pma_loss_of_signal_o;
    input usr_rx0_pma_pll_rst_n_i;
    input usr_rx0_rst_n_i;
    input [3:0] usr_rx0_test_i;
    output [7:0] usr_rx0_test_o;
    output usr_rx1_busy_o;
    input usr_rx1_ctrl_align_en_i;
    input usr_rx1_ctrl_align_sync_i;
    output [7:0] usr_rx1_ctrl_char_is_a_o;
    output usr_rx1_ctrl_char_is_aligned_o;
    output [7:0] usr_rx1_ctrl_char_is_comma_o;
    output [7:0] usr_rx1_ctrl_char_is_f_o;
    output [7:0] usr_rx1_ctrl_char_is_k_o;
    input usr_rx1_ctrl_dec_en_i;
    output [7:0] usr_rx1_ctrl_disp_err_o;
    input usr_rx1_ctrl_dscr_en_i;
    input usr_rx1_ctrl_el_buff_fifo_en_i;
    input usr_rx1_ctrl_el_buff_rst_i;
    output [7:0] usr_rx1_ctrl_not_in_table_o;
    input [1:0] usr_rx1_ctrl_ovs_bit_sel_i;
    input usr_rx1_ctrl_replace_en_i;
    output [63:0] usr_rx1_data_o;
    output usr_rx1_pll_lock_o;
    input usr_rx1_pma_cdr_rst_i;
    input usr_rx1_pma_ckgen_rst_n_i;
    output usr_rx1_pma_loss_of_signal_o;
    input usr_rx1_pma_pll_rst_n_i;
    input usr_rx1_rst_n_i;
    input [3:0] usr_rx1_test_i;
    output [7:0] usr_rx1_test_o;
    output usr_rx2_busy_o;
    input usr_rx2_ctrl_align_en_i;
    input usr_rx2_ctrl_align_sync_i;
    output [7:0] usr_rx2_ctrl_char_is_a_o;
    output usr_rx2_ctrl_char_is_aligned_o;
    output [7:0] usr_rx2_ctrl_char_is_comma_o;
    output [7:0] usr_rx2_ctrl_char_is_f_o;
    output [7:0] usr_rx2_ctrl_char_is_k_o;
    input usr_rx2_ctrl_dec_en_i;
    output [7:0] usr_rx2_ctrl_disp_err_o;
    input usr_rx2_ctrl_dscr_en_i;
    input usr_rx2_ctrl_el_buff_fifo_en_i;
    input usr_rx2_ctrl_el_buff_rst_i;
    output [7:0] usr_rx2_ctrl_not_in_table_o;
    input [1:0] usr_rx2_ctrl_ovs_bit_sel_i;
    input usr_rx2_ctrl_replace_en_i;
    output [63:0] usr_rx2_data_o;
    output usr_rx2_pll_lock_o;
    input usr_rx2_pma_cdr_rst_i;
    input usr_rx2_pma_ckgen_rst_n_i;
    output usr_rx2_pma_loss_of_signal_o;
    input usr_rx2_pma_pll_rst_n_i;
    input usr_rx2_rst_n_i;
    input [3:0] usr_rx2_test_i;
    output [7:0] usr_rx2_test_o;
    output usr_rx3_busy_o;
    input usr_rx3_ctrl_align_en_i;
    input usr_rx3_ctrl_align_sync_i;
    output [7:0] usr_rx3_ctrl_char_is_a_o;
    output usr_rx3_ctrl_char_is_aligned_o;
    output [7:0] usr_rx3_ctrl_char_is_comma_o;
    output [7:0] usr_rx3_ctrl_char_is_f_o;
    output [7:0] usr_rx3_ctrl_char_is_k_o;
    input usr_rx3_ctrl_dec_en_i;
    output [7:0] usr_rx3_ctrl_disp_err_o;
    input usr_rx3_ctrl_dscr_en_i;
    input usr_rx3_ctrl_el_buff_fifo_en_i;
    input usr_rx3_ctrl_el_buff_rst_i;
    output [7:0] usr_rx3_ctrl_not_in_table_o;
    input [1:0] usr_rx3_ctrl_ovs_bit_sel_i;
    input usr_rx3_ctrl_replace_en_i;
    output [63:0] usr_rx3_data_o;
    output usr_rx3_pll_lock_o;
    input usr_rx3_pma_cdr_rst_i;
    input usr_rx3_pma_ckgen_rst_n_i;
    output usr_rx3_pma_loss_of_signal_o;
    input usr_rx3_pma_pll_rst_n_i;
    input usr_rx3_rst_n_i;
    input [3:0] usr_rx3_test_i;
    output [7:0] usr_rx3_test_o;
    output usr_rx4_busy_o;
    input usr_rx4_ctrl_align_en_i;
    input usr_rx4_ctrl_align_sync_i;
    output [7:0] usr_rx4_ctrl_char_is_a_o;
    output usr_rx4_ctrl_char_is_aligned_o;
    output [7:0] usr_rx4_ctrl_char_is_comma_o;
    output [7:0] usr_rx4_ctrl_char_is_f_o;
    output [7:0] usr_rx4_ctrl_char_is_k_o;
    input usr_rx4_ctrl_dec_en_i;
    output [7:0] usr_rx4_ctrl_disp_err_o;
    input usr_rx4_ctrl_dscr_en_i;
    input usr_rx4_ctrl_el_buff_fifo_en_i;
    input usr_rx4_ctrl_el_buff_rst_i;
    output [7:0] usr_rx4_ctrl_not_in_table_o;
    input [1:0] usr_rx4_ctrl_ovs_bit_sel_i;
    input usr_rx4_ctrl_replace_en_i;
    output [63:0] usr_rx4_data_o;
    output usr_rx4_pll_lock_o;
    input usr_rx4_pma_cdr_rst_i;
    input usr_rx4_pma_ckgen_rst_n_i;
    output usr_rx4_pma_loss_of_signal_o;
    input usr_rx4_pma_pll_rst_n_i;
    input usr_rx4_rst_n_i;
    input [3:0] usr_rx4_test_i;
    output [7:0] usr_rx4_test_o;
    output usr_rx5_busy_o;
    input usr_rx5_ctrl_align_en_i;
    input usr_rx5_ctrl_align_sync_i;
    output [7:0] usr_rx5_ctrl_char_is_a_o;
    output usr_rx5_ctrl_char_is_aligned_o;
    output [7:0] usr_rx5_ctrl_char_is_comma_o;
    output [7:0] usr_rx5_ctrl_char_is_f_o;
    output [7:0] usr_rx5_ctrl_char_is_k_o;
    input usr_rx5_ctrl_dec_en_i;
    output [7:0] usr_rx5_ctrl_disp_err_o;
    input usr_rx5_ctrl_dscr_en_i;
    input usr_rx5_ctrl_el_buff_fifo_en_i;
    input usr_rx5_ctrl_el_buff_rst_i;
    output [7:0] usr_rx5_ctrl_not_in_table_o;
    input [1:0] usr_rx5_ctrl_ovs_bit_sel_i;
    input usr_rx5_ctrl_replace_en_i;
    output [63:0] usr_rx5_data_o;
    output usr_rx5_pll_lock_o;
    input usr_rx5_pma_cdr_rst_i;
    input usr_rx5_pma_ckgen_rst_n_i;
    output usr_rx5_pma_loss_of_signal_o;
    input usr_rx5_pma_pll_rst_n_i;
    input usr_rx5_rst_n_i;
    input [3:0] usr_rx5_test_i;
    output [7:0] usr_rx5_test_o;
    output usr_tx0_busy_o;
    input [7:0] usr_tx0_ctrl_char_is_k_i;
    input [7:0] usr_tx0_ctrl_enc_en_i;
    input [7:0] usr_tx0_ctrl_end_of_frame_i;
    input [7:0] usr_tx0_ctrl_end_of_multiframe_i;
    input usr_tx0_ctrl_replace_en_i;
    input [7:0] usr_tx0_ctrl_scr_en_i;
    input [63:0] usr_tx0_data_i;
    input usr_tx0_pma_clk_en_i;
    input usr_tx0_rst_n_i;
    input [3:0] usr_tx0_test_i;
    output [3:0] usr_tx0_test_o;
    output usr_tx1_busy_o;
    input [7:0] usr_tx1_ctrl_char_is_k_i;
    input [7:0] usr_tx1_ctrl_enc_en_i;
    input [7:0] usr_tx1_ctrl_end_of_frame_i;
    input [7:0] usr_tx1_ctrl_end_of_multiframe_i;
    input usr_tx1_ctrl_replace_en_i;
    input [7:0] usr_tx1_ctrl_scr_en_i;
    input [63:0] usr_tx1_data_i;
    input usr_tx1_pma_clk_en_i;
    input usr_tx1_rst_n_i;
    input [3:0] usr_tx1_test_i;
    output [3:0] usr_tx1_test_o;
    output usr_tx2_busy_o;
    input [7:0] usr_tx2_ctrl_char_is_k_i;
    input [7:0] usr_tx2_ctrl_enc_en_i;
    input [7:0] usr_tx2_ctrl_end_of_frame_i;
    input [7:0] usr_tx2_ctrl_end_of_multiframe_i;
    input usr_tx2_ctrl_replace_en_i;
    input [7:0] usr_tx2_ctrl_scr_en_i;
    input [63:0] usr_tx2_data_i;
    input usr_tx2_pma_clk_en_i;
    input usr_tx2_rst_n_i;
    input [3:0] usr_tx2_test_i;
    output [3:0] usr_tx2_test_o;
    output usr_tx3_busy_o;
    input [7:0] usr_tx3_ctrl_char_is_k_i;
    input [7:0] usr_tx3_ctrl_enc_en_i;
    input [7:0] usr_tx3_ctrl_end_of_frame_i;
    input [7:0] usr_tx3_ctrl_end_of_multiframe_i;
    input usr_tx3_ctrl_replace_en_i;
    input [7:0] usr_tx3_ctrl_scr_en_i;
    input [63:0] usr_tx3_data_i;
    input usr_tx3_pma_clk_en_i;
    input usr_tx3_rst_n_i;
    input [3:0] usr_tx3_test_i;
    output [3:0] usr_tx3_test_o;
    output usr_tx4_busy_o;
    input [7:0] usr_tx4_ctrl_char_is_k_i;
    input [7:0] usr_tx4_ctrl_enc_en_i;
    input [7:0] usr_tx4_ctrl_end_of_frame_i;
    input [7:0] usr_tx4_ctrl_end_of_multiframe_i;
    input usr_tx4_ctrl_replace_en_i;
    input [7:0] usr_tx4_ctrl_scr_en_i;
    input [63:0] usr_tx4_data_i;
    input usr_tx4_pma_clk_en_i;
    input usr_tx4_rst_n_i;
    input [3:0] usr_tx4_test_i;
    output [3:0] usr_tx4_test_o;
    output usr_tx5_busy_o;
    input [7:0] usr_tx5_ctrl_char_is_k_i;
    input [7:0] usr_tx5_ctrl_enc_en_i;
    input [7:0] usr_tx5_ctrl_end_of_frame_i;
    input [7:0] usr_tx5_ctrl_end_of_multiframe_i;
    input usr_tx5_ctrl_replace_en_i;
    input [7:0] usr_tx5_ctrl_scr_en_i;
    input [63:0] usr_tx5_data_i;
    input usr_tx5_pma_clk_en_i;
    input usr_tx5_rst_n_i;
    input [3:0] usr_tx5_test_i;
    output [3:0] usr_tx5_test_o;
    parameter cfg_main_i = 34'b0000000000000000000000000000000000;
    parameter cfg_rx0_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx1_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx2_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx3_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx4_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx5_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_tx0_i = 0;
    parameter cfg_tx1_i = 0;
    parameter cfg_tx2_i = 0;
    parameter cfg_tx3_i = 0;
    parameter cfg_tx4_i = 0;
    parameter cfg_tx5_i = 0;
    parameter location = "";
endmodule

(* blackbox *)
module NX_HSSL_U_FULL(hssl_clk_user_tx_i, hssl_clk_user_rx_i, hssl_clk_ref_i, hssl_clock_o, hssl_rclock_o, usr_dyn_cfg_en_i, usr_dyn_cfg_calibration_cs_n_i, usr_dyn_cfg_we_n_i, usr_dyn_cfg_wdata_sel_i, usr_pll_pma_rst_n_i, usr_pll_pma_pwr_down_n_i, usr_main_rst_n_i, usr_pll_lock_o, usr_pll_pma_lock_analog_o, usr_pll_ckfb_lock_o, usr_calibrate_pma_out_o, usr_main_async_debug_ack_i, usr_main_async_debug_req_o, scan_en_i, usr_tx0_ctrl_replace_en_i, usr_tx0_rst_n_i
, usr_tx0_busy_o, usr_tx0_ctrl_invalid_k_o, usr_tx0_ctrl_driver_pwrdwn_n_i, usr_tx0_pma_clk_en_i, usr_tx0_pma_tx_clk_o, usr_rx0_ctrl_dscr_en_i, usr_rx0_ctrl_dec_en_i, usr_rx0_ctrl_align_en_i, usr_rx0_ctrl_align_sync_i, usr_rx0_ctrl_replace_en_i, usr_rx0_ctrl_el_buff_rst_i, usr_rx0_rst_n_i, usr_rx0_pma_rst_n_i, usr_rx0_pma_m_eye_rst_i, usr_rx0_pma_pwr_down_n_i, usr_rx0_ctrl_char_is_aligned_o, usr_rx0_ctrl_valid_realign_o, usr_rx0_busy_o, usr_rx0_pma_loss_of_signal_o, usr_rx0_pma_ll_fast_locked_o, usr_rx0_pma_ll_slow_locked_o
, usr_rx0_pma_pll_lock_o, usr_rx0_pma_pll_lock_track_o, usr_tx1_ctrl_replace_en_i, usr_tx1_rst_n_i, usr_tx1_busy_o, usr_tx1_ctrl_invalid_k_o, usr_tx1_ctrl_driver_pwrdwn_n_i, usr_tx1_pma_clk_en_i, usr_tx1_pma_tx_clk_o, usr_rx1_ctrl_dscr_en_i, usr_rx1_ctrl_dec_en_i, usr_rx1_ctrl_align_en_i, usr_rx1_ctrl_align_sync_i, usr_rx1_ctrl_replace_en_i, usr_rx1_ctrl_el_buff_rst_i, usr_rx1_rst_n_i, usr_rx1_pma_rst_n_i, usr_rx1_pma_m_eye_rst_i, usr_rx1_pma_pwr_down_n_i, usr_rx1_ctrl_char_is_aligned_o, usr_rx1_ctrl_valid_realign_o
, usr_rx1_busy_o, usr_rx1_pma_loss_of_signal_o, usr_rx1_pma_ll_fast_locked_o, usr_rx1_pma_ll_slow_locked_o, usr_rx1_pma_pll_lock_o, usr_rx1_pma_pll_lock_track_o, usr_tx2_ctrl_replace_en_i, usr_tx2_rst_n_i, usr_tx2_busy_o, usr_tx2_ctrl_invalid_k_o, usr_tx2_ctrl_driver_pwrdwn_n_i, usr_tx2_pma_clk_en_i, usr_tx2_pma_tx_clk_o, usr_rx2_ctrl_dscr_en_i, usr_rx2_ctrl_dec_en_i, usr_rx2_ctrl_align_en_i, usr_rx2_ctrl_align_sync_i, usr_rx2_ctrl_replace_en_i, usr_rx2_ctrl_el_buff_rst_i, usr_rx2_rst_n_i, usr_rx2_pma_rst_n_i
, usr_rx2_pma_m_eye_rst_i, usr_rx2_pma_pwr_down_n_i, usr_rx2_ctrl_char_is_aligned_o, usr_rx2_ctrl_valid_realign_o, usr_rx2_busy_o, usr_rx2_pma_loss_of_signal_o, usr_rx2_pma_ll_fast_locked_o, usr_rx2_pma_ll_slow_locked_o, usr_rx2_pma_pll_lock_o, usr_rx2_pma_pll_lock_track_o, usr_tx3_ctrl_replace_en_i, usr_tx3_rst_n_i, usr_tx3_busy_o, usr_tx3_ctrl_invalid_k_o, usr_tx3_ctrl_driver_pwrdwn_n_i, usr_tx3_pma_clk_en_i, usr_tx3_pma_tx_clk_o, usr_rx3_ctrl_dscr_en_i, usr_rx3_ctrl_dec_en_i, usr_rx3_ctrl_align_en_i, usr_rx3_ctrl_align_sync_i
, usr_rx3_ctrl_replace_en_i, usr_rx3_ctrl_el_buff_rst_i, usr_rx3_rst_n_i, usr_rx3_pma_rst_n_i, usr_rx3_pma_m_eye_rst_i, usr_rx3_pma_pwr_down_n_i, usr_rx3_ctrl_char_is_aligned_o, usr_rx3_ctrl_valid_realign_o, usr_rx3_busy_o, usr_rx3_pma_loss_of_signal_o, usr_rx3_pma_ll_fast_locked_o, usr_rx3_pma_ll_slow_locked_o, usr_rx3_pma_pll_lock_o, usr_rx3_pma_pll_lock_track_o, usr_tx0_ctrl_enc_en_i, usr_tx0_ctrl_char_is_k_i, usr_tx0_ctrl_scr_en_i, usr_tx0_ctrl_end_of_multiframe_i, usr_tx0_ctrl_end_of_frame_i, usr_tx0_data_i, usr_rx0_data_o
, usr_rx0_ctrl_ovs_bit_sel_i, usr_rx0_ctrl_char_is_comma_o, usr_rx0_ctrl_char_is_k_o, usr_rx0_ctrl_not_in_table_o, usr_rx0_ctrl_disp_err_o, usr_rx0_ctrl_char_is_a_o, usr_rx0_ctrl_char_is_f_o, usr_rx0_test_o, usr_tx1_ctrl_enc_en_i, usr_tx1_ctrl_char_is_k_i, usr_tx1_ctrl_scr_en_i, usr_tx1_ctrl_end_of_multiframe_i, usr_tx1_ctrl_end_of_frame_i, usr_tx1_data_i, usr_rx1_data_o, usr_rx1_ctrl_ovs_bit_sel_i, usr_rx1_ctrl_char_is_comma_o, usr_rx1_ctrl_char_is_k_o, usr_rx1_ctrl_not_in_table_o, usr_rx1_ctrl_disp_err_o, usr_rx1_ctrl_char_is_a_o
, usr_rx1_ctrl_char_is_f_o, usr_rx1_test_o, usr_tx2_ctrl_enc_en_i, usr_tx2_ctrl_char_is_k_i, usr_tx2_ctrl_scr_en_i, usr_tx2_ctrl_end_of_multiframe_i, usr_tx2_ctrl_end_of_frame_i, usr_tx2_data_i, usr_rx2_data_o, usr_rx2_ctrl_ovs_bit_sel_i, usr_rx2_ctrl_char_is_comma_o, usr_rx2_ctrl_char_is_k_o, usr_rx2_ctrl_not_in_table_o, usr_rx2_ctrl_disp_err_o, usr_rx2_ctrl_char_is_a_o, usr_rx2_ctrl_char_is_f_o, usr_rx2_test_o, usr_tx3_ctrl_enc_en_i, usr_tx3_ctrl_char_is_k_i, usr_tx3_ctrl_scr_en_i, usr_tx3_ctrl_end_of_multiframe_i
, usr_tx3_ctrl_end_of_frame_i, usr_tx3_data_i, usr_rx3_data_o, usr_rx3_ctrl_ovs_bit_sel_i, usr_rx3_ctrl_char_is_comma_o, usr_rx3_ctrl_char_is_k_o, usr_rx3_ctrl_not_in_table_o, usr_rx3_ctrl_disp_err_o, usr_rx3_ctrl_char_is_a_o, usr_rx3_ctrl_char_is_f_o, usr_rx3_test_o, usr_dyn_cfg_addr_i, usr_dyn_cfg_wdata_i, usr_main_async_debug_lane_sel_i, usr_main_rx_pma_ll_out_o, scan_in_i, scan_out_o, usr_rx0_ctrl_debug_sel_i, usr_rx1_ctrl_debug_sel_i, usr_rx2_ctrl_debug_sel_i, usr_rx3_ctrl_debug_sel_i
, usr_dyn_cfg_lane_cs_n_i);
    input hssl_clk_ref_i;
    input hssl_clk_user_rx_i;
    input hssl_clk_user_tx_i;
    output hssl_clock_o;
    output hssl_rclock_o;
    input scan_en_i;
    input [7:0] scan_in_i;
    output [7:0] scan_out_o;
    output usr_calibrate_pma_out_o;
    input [3:0] usr_dyn_cfg_addr_i;
    input usr_dyn_cfg_calibration_cs_n_i;
    input usr_dyn_cfg_en_i;
    input [3:0] usr_dyn_cfg_lane_cs_n_i;
    input [11:0] usr_dyn_cfg_wdata_i;
    input usr_dyn_cfg_wdata_sel_i;
    input usr_dyn_cfg_we_n_i;
    input usr_main_async_debug_ack_i;
    input [1:0] usr_main_async_debug_lane_sel_i;
    output usr_main_async_debug_req_o;
    input usr_main_rst_n_i;
    output [19:0] usr_main_rx_pma_ll_out_o;
    output usr_pll_ckfb_lock_o;
    output usr_pll_lock_o;
    output usr_pll_pma_lock_analog_o;
    input usr_pll_pma_pwr_down_n_i;
    input usr_pll_pma_rst_n_i;
    output usr_rx0_busy_o;
    input usr_rx0_ctrl_align_en_i;
    input usr_rx0_ctrl_align_sync_i;
    output [7:0] usr_rx0_ctrl_char_is_a_o;
    output usr_rx0_ctrl_char_is_aligned_o;
    output [7:0] usr_rx0_ctrl_char_is_comma_o;
    output [7:0] usr_rx0_ctrl_char_is_f_o;
    output [7:0] usr_rx0_ctrl_char_is_k_o;
    input [2:0] usr_rx0_ctrl_debug_sel_i;
    input usr_rx0_ctrl_dec_en_i;
    output [7:0] usr_rx0_ctrl_disp_err_o;
    input usr_rx0_ctrl_dscr_en_i;
    input usr_rx0_ctrl_el_buff_rst_i;
    output [7:0] usr_rx0_ctrl_not_in_table_o;
    input [1:0] usr_rx0_ctrl_ovs_bit_sel_i;
    input usr_rx0_ctrl_replace_en_i;
    output usr_rx0_ctrl_valid_realign_o;
    output [63:0] usr_rx0_data_o;
    output usr_rx0_pma_ll_fast_locked_o;
    output usr_rx0_pma_ll_slow_locked_o;
    output usr_rx0_pma_loss_of_signal_o;
    input usr_rx0_pma_m_eye_rst_i;
    output usr_rx0_pma_pll_lock_o;
    output usr_rx0_pma_pll_lock_track_o;
    input usr_rx0_pma_pwr_down_n_i;
    input usr_rx0_pma_rst_n_i;
    input usr_rx0_rst_n_i;
    output [7:0] usr_rx0_test_o;
    output usr_rx1_busy_o;
    input usr_rx1_ctrl_align_en_i;
    input usr_rx1_ctrl_align_sync_i;
    output [7:0] usr_rx1_ctrl_char_is_a_o;
    output usr_rx1_ctrl_char_is_aligned_o;
    output [7:0] usr_rx1_ctrl_char_is_comma_o;
    output [7:0] usr_rx1_ctrl_char_is_f_o;
    output [7:0] usr_rx1_ctrl_char_is_k_o;
    input [2:0] usr_rx1_ctrl_debug_sel_i;
    input usr_rx1_ctrl_dec_en_i;
    output [7:0] usr_rx1_ctrl_disp_err_o;
    input usr_rx1_ctrl_dscr_en_i;
    input usr_rx1_ctrl_el_buff_rst_i;
    output [7:0] usr_rx1_ctrl_not_in_table_o;
    input [1:0] usr_rx1_ctrl_ovs_bit_sel_i;
    input usr_rx1_ctrl_replace_en_i;
    output usr_rx1_ctrl_valid_realign_o;
    output [63:0] usr_rx1_data_o;
    output usr_rx1_pma_ll_fast_locked_o;
    output usr_rx1_pma_ll_slow_locked_o;
    output usr_rx1_pma_loss_of_signal_o;
    input usr_rx1_pma_m_eye_rst_i;
    output usr_rx1_pma_pll_lock_o;
    output usr_rx1_pma_pll_lock_track_o;
    input usr_rx1_pma_pwr_down_n_i;
    input usr_rx1_pma_rst_n_i;
    input usr_rx1_rst_n_i;
    output [7:0] usr_rx1_test_o;
    output usr_rx2_busy_o;
    input usr_rx2_ctrl_align_en_i;
    input usr_rx2_ctrl_align_sync_i;
    output [7:0] usr_rx2_ctrl_char_is_a_o;
    output usr_rx2_ctrl_char_is_aligned_o;
    output [7:0] usr_rx2_ctrl_char_is_comma_o;
    output [7:0] usr_rx2_ctrl_char_is_f_o;
    output [7:0] usr_rx2_ctrl_char_is_k_o;
    input [2:0] usr_rx2_ctrl_debug_sel_i;
    input usr_rx2_ctrl_dec_en_i;
    output [7:0] usr_rx2_ctrl_disp_err_o;
    input usr_rx2_ctrl_dscr_en_i;
    input usr_rx2_ctrl_el_buff_rst_i;
    output [7:0] usr_rx2_ctrl_not_in_table_o;
    input [1:0] usr_rx2_ctrl_ovs_bit_sel_i;
    input usr_rx2_ctrl_replace_en_i;
    output usr_rx2_ctrl_valid_realign_o;
    output [63:0] usr_rx2_data_o;
    output usr_rx2_pma_ll_fast_locked_o;
    output usr_rx2_pma_ll_slow_locked_o;
    output usr_rx2_pma_loss_of_signal_o;
    input usr_rx2_pma_m_eye_rst_i;
    output usr_rx2_pma_pll_lock_o;
    output usr_rx2_pma_pll_lock_track_o;
    input usr_rx2_pma_pwr_down_n_i;
    input usr_rx2_pma_rst_n_i;
    input usr_rx2_rst_n_i;
    output [7:0] usr_rx2_test_o;
    output usr_rx3_busy_o;
    input usr_rx3_ctrl_align_en_i;
    input usr_rx3_ctrl_align_sync_i;
    output [7:0] usr_rx3_ctrl_char_is_a_o;
    output usr_rx3_ctrl_char_is_aligned_o;
    output [7:0] usr_rx3_ctrl_char_is_comma_o;
    output [7:0] usr_rx3_ctrl_char_is_f_o;
    output [7:0] usr_rx3_ctrl_char_is_k_o;
    input [2:0] usr_rx3_ctrl_debug_sel_i;
    input usr_rx3_ctrl_dec_en_i;
    output [7:0] usr_rx3_ctrl_disp_err_o;
    input usr_rx3_ctrl_dscr_en_i;
    input usr_rx3_ctrl_el_buff_rst_i;
    output [7:0] usr_rx3_ctrl_not_in_table_o;
    input [1:0] usr_rx3_ctrl_ovs_bit_sel_i;
    input usr_rx3_ctrl_replace_en_i;
    output usr_rx3_ctrl_valid_realign_o;
    output [63:0] usr_rx3_data_o;
    output usr_rx3_pma_ll_fast_locked_o;
    output usr_rx3_pma_ll_slow_locked_o;
    output usr_rx3_pma_loss_of_signal_o;
    input usr_rx3_pma_m_eye_rst_i;
    output usr_rx3_pma_pll_lock_o;
    output usr_rx3_pma_pll_lock_track_o;
    input usr_rx3_pma_pwr_down_n_i;
    input usr_rx3_pma_rst_n_i;
    input usr_rx3_rst_n_i;
    output [7:0] usr_rx3_test_o;
    output usr_tx0_busy_o;
    input [7:0] usr_tx0_ctrl_char_is_k_i;
    input usr_tx0_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx0_ctrl_enc_en_i;
    input [7:0] usr_tx0_ctrl_end_of_frame_i;
    input [7:0] usr_tx0_ctrl_end_of_multiframe_i;
    output usr_tx0_ctrl_invalid_k_o;
    input usr_tx0_ctrl_replace_en_i;
    input [7:0] usr_tx0_ctrl_scr_en_i;
    input [63:0] usr_tx0_data_i;
    input usr_tx0_pma_clk_en_i;
    output usr_tx0_pma_tx_clk_o;
    input usr_tx0_rst_n_i;
    output usr_tx1_busy_o;
    input [7:0] usr_tx1_ctrl_char_is_k_i;
    input usr_tx1_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx1_ctrl_enc_en_i;
    input [7:0] usr_tx1_ctrl_end_of_frame_i;
    input [7:0] usr_tx1_ctrl_end_of_multiframe_i;
    output usr_tx1_ctrl_invalid_k_o;
    input usr_tx1_ctrl_replace_en_i;
    input [7:0] usr_tx1_ctrl_scr_en_i;
    input [63:0] usr_tx1_data_i;
    input usr_tx1_pma_clk_en_i;
    output usr_tx1_pma_tx_clk_o;
    input usr_tx1_rst_n_i;
    output usr_tx2_busy_o;
    input [7:0] usr_tx2_ctrl_char_is_k_i;
    input usr_tx2_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx2_ctrl_enc_en_i;
    input [7:0] usr_tx2_ctrl_end_of_frame_i;
    input [7:0] usr_tx2_ctrl_end_of_multiframe_i;
    output usr_tx2_ctrl_invalid_k_o;
    input usr_tx2_ctrl_replace_en_i;
    input [7:0] usr_tx2_ctrl_scr_en_i;
    input [63:0] usr_tx2_data_i;
    input usr_tx2_pma_clk_en_i;
    output usr_tx2_pma_tx_clk_o;
    input usr_tx2_rst_n_i;
    output usr_tx3_busy_o;
    input [7:0] usr_tx3_ctrl_char_is_k_i;
    input usr_tx3_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx3_ctrl_enc_en_i;
    input [7:0] usr_tx3_ctrl_end_of_frame_i;
    input [7:0] usr_tx3_ctrl_end_of_multiframe_i;
    output usr_tx3_ctrl_invalid_k_o;
    input usr_tx3_ctrl_replace_en_i;
    input [7:0] usr_tx3_ctrl_scr_en_i;
    input [63:0] usr_tx3_data_i;
    input usr_tx3_pma_clk_en_i;
    output usr_tx3_pma_tx_clk_o;
    input usr_tx3_rst_n_i;
    parameter cfg_dyn_all_rx_pma_m_eye_coarse_ena_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_dn_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_fine_ena_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_step_i = 4'b0000;
    parameter cfg_dyn_all_rx_pma_m_eye_up_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_threshold_1 = 5'b00000;
    parameter cfg_dyn_all_rx_pma_threshold_2 = 5'b00000;
    parameter cfg_dyn_all_rx_pma_trim_locked_i = 3'b000;
    parameter cfg_dyn_all_rx_pma_trim_mode_i = 2'b00;
    parameter cfg_dyn_all_rx_pma_trim_unlocked_i = 3'b000;
    parameter cfg_dyn_rx0_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx0_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx1_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx2_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx3_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_tx0_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx0_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx0_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx0_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx0_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx0_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx0_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx0_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx0_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx0_pma_pre_sign_i = 1'b0;
    parameter cfg_dyn_tx1_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx1_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx1_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx1_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx1_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx1_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx1_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx1_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx1_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx1_pma_pre_sign_i = 1'b0;
    parameter cfg_dyn_tx2_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx2_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx2_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx2_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx2_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx2_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx2_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx2_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx2_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx2_pma_pre_sign_i = 1'b0;
    parameter cfg_dyn_tx3_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx3_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx3_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx3_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx3_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx3_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx3_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx3_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx3_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx3_pma_pre_sign_i = 1'b0;
    parameter cfg_main_clk_to_fabric_div_en_i = 1'b0;
    parameter cfg_main_clk_to_fabric_div_mode_i = 1'b0;
    parameter cfg_main_clk_to_fabric_sel_i = 1'b0;
    parameter cfg_main_rclk_to_fabric_sel_i = 2'b00;
    parameter cfg_main_use_only_usr_clock_i = 1'b0;
    parameter cfg_pcs_ovs_en_i = 1'b0;
    parameter cfg_pcs_ovs_mode_i = 1'b0;
    parameter cfg_pcs_pll_lock_ppm_i = 3'b000;
    parameter cfg_pcs_word_len_i = 2'b00;
    parameter cfg_pll_pma_ckref_ext_i = 1'b0;
    parameter cfg_pll_pma_cpump_i = 4'b0000;
    parameter cfg_pll_pma_divl_i = 2'b00;
    parameter cfg_pll_pma_divm_i = 1'b0;
    parameter cfg_pll_pma_divn_i = 2'b00;
    parameter cfg_pll_pma_gbx_en_i = 1'b0;
    parameter cfg_pll_pma_int_data_len_i = 1'b0;
    parameter cfg_pll_pma_lvds_en_i = 1'b0;
    parameter cfg_pll_pma_lvds_mux_i = 1'b0;
    parameter cfg_pll_pma_mux_ckref_i = 1'b0;
    parameter cfg_rx0_gearbox_en_i = 1'b0;
    parameter cfg_rx0_gearbox_mode_i = 1'b0;
    parameter cfg_rx0_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx0_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx0_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx0_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx0_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx0_pcs_debug_en_i = 1'b0;
    parameter cfg_rx0_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx0_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx0_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx0_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx0_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx0_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx0_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx0_pcs_loopback_i = 1'b0;
    parameter cfg_rx0_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx0_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx0_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx0_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx0_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx0_pcs_polarity_i = 1'b0;
    parameter cfg_rx0_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx0_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx0_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx0_pma_clk_pos_i = 1'b0;
    parameter cfg_rx0_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx0_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx0_pma_dco_divl_i = 2'b00;
    parameter cfg_rx0_pma_dco_divm_i = 1'b0;
    parameter cfg_rx0_pma_dco_divn_i = 2'b00;
    parameter cfg_rx0_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx0_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx0_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx0_pma_loopback_i = 1'b0;
    parameter cfg_rx0_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx0_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx0_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx0_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx0_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx0_pma_pll_divf_i = 2'b00;
    parameter cfg_rx0_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx0_pma_pll_divm_i = 2'b00;
    parameter cfg_rx0_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx0_pma_pll_divn_i = 1'b0;
    parameter cfg_rx1_gearbox_en_i = 1'b0;
    parameter cfg_rx1_gearbox_mode_i = 1'b0;
    parameter cfg_rx1_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx1_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx1_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx1_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx1_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx1_pcs_debug_en_i = 1'b0;
    parameter cfg_rx1_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx1_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx1_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx1_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx1_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx1_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx1_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx1_pcs_loopback_i = 1'b0;
    parameter cfg_rx1_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx1_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx1_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx1_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx1_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx1_pcs_polarity_i = 1'b0;
    parameter cfg_rx1_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx1_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx1_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx1_pma_clk_pos_i = 1'b0;
    parameter cfg_rx1_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx1_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx1_pma_dco_divl_i = 2'b00;
    parameter cfg_rx1_pma_dco_divm_i = 1'b0;
    parameter cfg_rx1_pma_dco_divn_i = 2'b00;
    parameter cfg_rx1_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx1_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx1_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx1_pma_loopback_i = 1'b0;
    parameter cfg_rx1_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx1_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx1_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx1_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx1_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx1_pma_pll_divf_i = 2'b00;
    parameter cfg_rx1_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx1_pma_pll_divm_i = 2'b00;
    parameter cfg_rx1_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx1_pma_pll_divn_i = 1'b0;
    parameter cfg_rx2_gearbox_en_i = 1'b0;
    parameter cfg_rx2_gearbox_mode_i = 1'b0;
    parameter cfg_rx2_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx2_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx2_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx2_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx2_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx2_pcs_debug_en_i = 1'b0;
    parameter cfg_rx2_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx2_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx2_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx2_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx2_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx2_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx2_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx2_pcs_loopback_i = 1'b0;
    parameter cfg_rx2_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx2_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx2_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx2_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx2_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx2_pcs_polarity_i = 1'b0;
    parameter cfg_rx2_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx2_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx2_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx2_pma_clk_pos_i = 1'b0;
    parameter cfg_rx2_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx2_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx2_pma_dco_divl_i = 2'b00;
    parameter cfg_rx2_pma_dco_divm_i = 1'b0;
    parameter cfg_rx2_pma_dco_divn_i = 2'b00;
    parameter cfg_rx2_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx2_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx2_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx2_pma_loopback_i = 1'b0;
    parameter cfg_rx2_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx2_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx2_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx2_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx2_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx2_pma_pll_divf_i = 2'b00;
    parameter cfg_rx2_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx2_pma_pll_divm_i = 2'b00;
    parameter cfg_rx2_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx2_pma_pll_divn_i = 1'b0;
    parameter cfg_rx3_gearbox_en_i = 1'b0;
    parameter cfg_rx3_gearbox_mode_i = 1'b0;
    parameter cfg_rx3_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx3_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx3_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx3_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx3_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx3_pcs_debug_en_i = 1'b0;
    parameter cfg_rx3_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx3_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx3_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx3_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx3_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx3_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx3_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx3_pcs_loopback_i = 1'b0;
    parameter cfg_rx3_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx3_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx3_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx3_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx3_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx3_pcs_polarity_i = 1'b0;
    parameter cfg_rx3_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx3_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx3_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx3_pma_clk_pos_i = 1'b0;
    parameter cfg_rx3_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx3_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx3_pma_dco_divl_i = 2'b00;
    parameter cfg_rx3_pma_dco_divm_i = 1'b0;
    parameter cfg_rx3_pma_dco_divn_i = 2'b00;
    parameter cfg_rx3_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx3_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx3_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx3_pma_loopback_i = 1'b0;
    parameter cfg_rx3_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx3_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx3_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx3_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx3_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx3_pma_pll_divf_i = 2'b00;
    parameter cfg_rx3_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx3_pma_pll_divm_i = 2'b00;
    parameter cfg_rx3_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx3_pma_pll_divn_i = 1'b0;
    parameter cfg_test_mode_i = 2'b00;
    parameter cfg_tx0_gearbox_en_i = 1'b0;
    parameter cfg_tx0_gearbox_mode_i = 1'b0;
    parameter cfg_tx0_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx0_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx0_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx0_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx0_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx0_pcs_loopback_i = 1'b0;
    parameter cfg_tx0_pcs_polarity_i = 1'b0;
    parameter cfg_tx0_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx0_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx0_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx0_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx0_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx0_pma_clk_pos_i = 1'b0;
    parameter cfg_tx0_pma_loopback_i = 1'b0;
    parameter cfg_tx1_gearbox_en_i = 1'b0;
    parameter cfg_tx1_gearbox_mode_i = 1'b0;
    parameter cfg_tx1_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx1_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx1_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx1_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx1_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx1_pcs_loopback_i = 1'b0;
    parameter cfg_tx1_pcs_polarity_i = 1'b0;
    parameter cfg_tx1_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx1_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx1_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx1_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx1_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx1_pma_clk_pos_i = 1'b0;
    parameter cfg_tx1_pma_loopback_i = 1'b0;
    parameter cfg_tx2_gearbox_en_i = 1'b0;
    parameter cfg_tx2_gearbox_mode_i = 1'b0;
    parameter cfg_tx2_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx2_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx2_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx2_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx2_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx2_pcs_loopback_i = 1'b0;
    parameter cfg_tx2_pcs_polarity_i = 1'b0;
    parameter cfg_tx2_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx2_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx2_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx2_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx2_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx2_pma_clk_pos_i = 1'b0;
    parameter cfg_tx2_pma_loopback_i = 1'b0;
    parameter cfg_tx3_gearbox_en_i = 1'b0;
    parameter cfg_tx3_gearbox_mode_i = 1'b0;
    parameter cfg_tx3_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx3_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx3_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx3_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx3_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx3_pcs_loopback_i = 1'b0;
    parameter cfg_tx3_pcs_polarity_i = 1'b0;
    parameter cfg_tx3_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx3_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx3_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx3_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx3_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx3_pma_clk_pos_i = 1'b0;
    parameter cfg_tx3_pma_loopback_i = 1'b0;
    parameter location = "";
    parameter rx_usrclk_use_pcs_clk_2 = 1'b0;
    parameter tx_usrclk_use_pcs_clk_2 = 1'b0;
endmodule

(* blackbox *)
module NX_IOB(I, C, T, O, IO);
    input C;
    input I;
    inout IO;
    output O;
    input T;
    parameter differential = "";
    parameter drive = "";
    parameter dynDrive = "";
    parameter dynInput = "";
    parameter dynTerm = "";
    parameter extra = 3;
    parameter inputDelayLine = "";
    parameter inputDelayOn = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter outputDelayOn = "";
    parameter slewRate = "";
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_IOB_I(C, T, IO, O);
    input C;
    input IO;
    output O;
    input T;
    parameter differential = "";
    parameter drive = "";
    parameter dynDrive = "";
    parameter dynInput = "";
    parameter dynTerm = "";
    parameter extra = 1;
    parameter inputDelayLine = "";
    parameter inputDelayOn = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter outputDelayOn = "";
    parameter slewRate = "";
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_IOB_O(I, C, T, IO);
    input C;
    input I;
    output IO;
    input T;
    parameter differential = "";
    parameter drive = "";
    parameter dynDrive = "";
    parameter dynInput = "";
    parameter dynTerm = "";
    parameter extra = 2;
    parameter inputDelayLine = "";
    parameter inputDelayOn = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter outputDelayOn = "";
    parameter slewRate = "";
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_IOM_BIN2GRP(GS, DS, GVON, GVIN, GVDN, PA, LA);
    input [1:0] DS;
    input GS;
    output [2:0] GVDN;
    output [2:0] GVIN;
    output [2:0] GVON;
    input [5:0] LA;
    output [3:0] PA;
endmodule

(* blackbox *)
module NX_IOM_CONTROL(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1, C2RW2, C2RW3
, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, CCK, DCK, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, SPI1, SPI2, SPI3, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1
, DRO2, DRO3, DRO4, DRO5, DRO6, CAL, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16
, LINK17, LINK18, LINK19, LINK20, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input SPI1;
    input SPI2;
    input SPI3;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter inv_di_fclk1 = 1'b0;
    parameter inv_di_fclk2 = 1'b0;
    parameter latency1 = 1'b0;
    parameter latency2 = 1'b0;
    parameter location = "";
    parameter mode_cpath = "";
    parameter mode_epath = "";
    parameter mode_io_cal = 1'b0;
    parameter mode_rpath = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_tpath = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_CONTROL_L(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1, C2RW2, C2RW3
, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, CCK, DCK, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1, DRO2, DRO3, DRO4
, DRO5, DRO6, CAL, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16, LINK17, LINK18, LINK19
, LINK20, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter inv_di_fclk1 = 1'b0;
    parameter inv_di_fclk2 = 1'b0;
    parameter latency1 = 1'b0;
    parameter latency2 = 1'b0;
    parameter location = "";
    parameter mode_cpath = "";
    parameter mode_epath = "";
    parameter mode_io_cal = 1'b0;
    parameter mode_rpath = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_tpath = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_CONTROL_M(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1, C2RW2, C2RW3
, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, CCK, DCK, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, SPI1, SPI2, SPI3, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1
, DRO2, DRO3, DRO4, DRO5, DRO6, CAL, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16
, LINK17, LINK18, LINK19, LINK20, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input SPI1;
    input SPI2;
    input SPI3;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter inv_di_fclk1 = 1'b0;
    parameter inv_di_fclk2 = 1'b0;
    parameter latency1 = 1'b0;
    parameter latency2 = 1'b0;
    parameter location = "";
    parameter mode_cpath = "";
    parameter mode_epath = "";
    parameter mode_io_cal = 1'b0;
    parameter mode_rpath = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_tpath = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_CONTROL_U(ALCK1, ALCK2, ALCK3, LDSCK1, LDSCK2, LDSCK3, SWRX1CK, SWRX2CK, FCK1, FCK2, FDCK, CCK, DQ1CI1, DQ1CI2, DQ1CI3, DQ1CI4, DQ1CI5, DQ1CI6, DQ1CI7, DQ1CI8, DQ2CI1
, DQ2CI2, DQ2CI3, DQ2CI4, DQ2CI5, DQ2CI6, DQ2CI7, DQ2CI8, DQ3CI1, DQ3CI2, DQ3CI3, DQ3CI4, DQ3CI5, DQ3CI6, DQ3CI7, DQ3CI8, DQS1CI1, DQS1CI2, DQS1CI3, DQS1CI4, DQS1CI5, DQS1CI6
, DQS1CI7, DQS1CI8, DQS2CI1, DQS2CI2, DQS2CI3, DQS2CI4, DQS2CI5, DQS2CI6, DQS2CI7, DQS2CI8, DQS3CI1, DQS3CI2, DQS3CI3, DQS3CI4, DQS3CI5, DQS3CI6, DQS3CI7, DQS3CI8, LD1RN, LD2RN, LD3RN
, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DCRN, LE, SE, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3, DRA4, DRO1CSN
, DRO2CSN, DRO3CSN, DRI1CSN, DRI2CSN, DRI3CSN, DRDPA1CSN, DRDPA2CSN, DRDPA3CSN, DRCCSN, DRWDS, DRWEN, DRE, CA1P1, CA1P2, CA1P3, CA1P4, CA2P1, CA2P2, CA2P3, CA2P4, CA1N1
, CA1N2, CA1N3, CA1N4, CA2N1, CA2N2, CA2N3, CA2N4, CA1T1, CA1T2, CA1T3, CA1T4, CA2T1, CA2T2, CA2T3, CA2T4, CA1D1, CA1D2, CA1D3, CA1D4, CA1D5, CA1D6
, CA2D1, CA2D2, CA2D3, CA2D4, CA2D5, CA2D6, CKO1, CKO2, FLD, FLG, AL1D, AL2D, AL3D, AL1T, AL2T, AL3T, DCL, DRO1, DRO2, DRO3, DRO4
, DRO5, DRO6, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16, LINK17, LINK18, LINK19, LINK20
, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output AL1D;
    output AL1T;
    output AL2D;
    output AL2T;
    output AL3D;
    output AL3T;
    input ALCK1;
    input ALCK2;
    input ALCK3;
    input CA1D1;
    input CA1D2;
    input CA1D3;
    input CA1D4;
    input CA1D5;
    input CA1D6;
    input CA1N1;
    input CA1N2;
    input CA1N3;
    input CA1N4;
    input CA1P1;
    input CA1P2;
    input CA1P3;
    input CA1P4;
    input CA1T1;
    input CA1T2;
    input CA1T3;
    input CA1T4;
    input CA2D1;
    input CA2D2;
    input CA2D3;
    input CA2D4;
    input CA2D5;
    input CA2D6;
    input CA2N1;
    input CA2N2;
    input CA2N3;
    input CA2N4;
    input CA2P1;
    input CA2P2;
    input CA2P3;
    input CA2P4;
    input CA2T1;
    input CA2T2;
    input CA2T3;
    input CA2T4;
    input CCK;
    output CKO1;
    output CKO2;
    output DCL;
    input DCRN;
    input DQ1CI1;
    input DQ1CI2;
    input DQ1CI3;
    input DQ1CI4;
    input DQ1CI5;
    input DQ1CI6;
    input DQ1CI7;
    input DQ1CI8;
    input DQ2CI1;
    input DQ2CI2;
    input DQ2CI3;
    input DQ2CI4;
    input DQ2CI5;
    input DQ2CI6;
    input DQ2CI7;
    input DQ2CI8;
    input DQ3CI1;
    input DQ3CI2;
    input DQ3CI3;
    input DQ3CI4;
    input DQ3CI5;
    input DQ3CI6;
    input DQ3CI7;
    input DQ3CI8;
    input DQS1CI1;
    input DQS1CI2;
    input DQS1CI3;
    input DQS1CI4;
    input DQS1CI5;
    input DQS1CI6;
    input DQS1CI7;
    input DQS1CI8;
    input DQS2CI1;
    input DQS2CI2;
    input DQS2CI3;
    input DQS2CI4;
    input DQS2CI5;
    input DQS2CI6;
    input DQS2CI7;
    input DQS2CI8;
    input DQS3CI1;
    input DQS3CI2;
    input DQS3CI3;
    input DQS3CI4;
    input DQS3CI5;
    input DQS3CI6;
    input DQS3CI7;
    input DQS3CI8;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRCCSN;
    input DRDPA1CSN;
    input DRDPA2CSN;
    input DRDPA3CSN;
    input DRE;
    input DRI1;
    input DRI1CSN;
    input DRI2;
    input DRI2CSN;
    input DRI3;
    input DRI3CSN;
    input DRI4;
    input DRI5;
    input DRI6;
    output DRO1;
    input DRO1CSN;
    output DRO2;
    input DRO2CSN;
    output DRO3;
    input DRO3CSN;
    output DRO4;
    output DRO5;
    output DRO6;
    input DRWDS;
    input DRWEN;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    input FCK1;
    input FCK2;
    input FDCK;
    output FLD;
    output FLG;
    input FZ;
    input LD1RN;
    input LD2RN;
    input LD3RN;
    input LDSCK1;
    input LDSCK2;
    input LDSCK3;
    input LE;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input SE;
    input SWRX1CK;
    input SWRX2CK;
    parameter cal_delay1 = "";
    parameter cal_delay2 = "";
    parameter div1 = 3'b000;
    parameter div2 = 3'b000;
    parameter div3 = 3'b000;
    parameter div_swrx1 = 3'b000;
    parameter div_swrx2 = 3'b000;
    parameter inv_ld_sck1 = 1'b0;
    parameter inv_ld_sck2 = 1'b0;
    parameter inv_ld_sck3 = 1'b0;
    parameter link_ld_12 = 1'b0;
    parameter link_ld_23 = 1'b0;
    parameter location = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_side3 = 0;
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_dc_clk = 2'b00;
    parameter sel_ld_fck1 = 2'b00;
    parameter sel_ld_fck2 = 2'b00;
    parameter sel_ld_fck3 = 2'b00;
    parameter sel_sw_fck1 = 2'b00;
    parameter sel_sw_fck2 = 2'b00;
    parameter use_dc = 1'b0;
endmodule

(* blackbox *)
module NX_IOM_DRIVER(EI1, EI2, EI3, EI4, EI5, EL, ER, CI1, CI2, CI3, CI4, CI5, CL, CR, CTI, RI, RL, RR, CO, EO, RO1
, RO2, RO3, RO4, RO5, CTO, LINK);
    input CI1;
    input CI2;
    input CI3;
    input CI4;
    input CI5;
    input CL;
    output CO;
    input CR;
    input CTI;
    output CTO;
    input EI1;
    input EI2;
    input EI3;
    input EI4;
    input EI5;
    input EL;
    output EO;
    input ER;
    inout [41:0] LINK;
    input RI;
    input RL;
    output RO1;
    output RO2;
    output RO3;
    output RO4;
    output RO5;
    input RR;
    parameter chained = 1'b0;
    parameter cpath_edge = 1'b0;
    parameter cpath_init = 1'b0;
    parameter cpath_inv = 1'b0;
    parameter cpath_load = 1'b0;
    parameter cpath_mode = 4'b0000;
    parameter cpath_sync = 1'b0;
    parameter epath_dynamic = 1'b0;
    parameter epath_edge = 1'b0;
    parameter epath_init = 1'b0;
    parameter epath_load = 1'b0;
    parameter epath_mode = 4'b0000;
    parameter epath_sync = 1'b0;
    parameter location = "";
    parameter rpath_dynamic = 1'b0;
    parameter rpath_edge = 1'b0;
    parameter rpath_init = 1'b0;
    parameter rpath_load = 1'b0;
    parameter rpath_mode = 4'b0000;
    parameter rpath_sync = 1'b0;
    parameter symbol = "";
    parameter tpath_mode = 2'b00;
    parameter variant = "";
endmodule

(* blackbox *)
module NX_IOM_DRIVER_M(EI1, EI2, EI3, EI4, EI5, EL, ER, CI1, CI2, CI3, CI4, CI5, CL, CR, CTI, RI, RL, RR, CO, EO, RO1
, RO2, RO3, RO4, RO5, CTO, LINK);
    input CI1;
    input CI2;
    input CI3;
    input CI4;
    input CI5;
    input CL;
    output CO;
    input CR;
    input CTI;
    output CTO;
    input EI1;
    input EI2;
    input EI3;
    input EI4;
    input EI5;
    input EL;
    output EO;
    input ER;
    inout [41:0] LINK;
    input RI;
    input RL;
    output RO1;
    output RO2;
    output RO3;
    output RO4;
    output RO5;
    input RR;
    parameter chained = 1'b0;
    parameter cpath_edge = 1'b0;
    parameter cpath_init = 1'b0;
    parameter cpath_inv = 1'b0;
    parameter cpath_load = 1'b0;
    parameter cpath_mode = 4'b0000;
    parameter cpath_sync = 1'b0;
    parameter epath_dynamic = 1'b0;
    parameter epath_edge = 1'b0;
    parameter epath_init = 1'b0;
    parameter epath_load = 1'b0;
    parameter epath_mode = 4'b0000;
    parameter epath_sync = 1'b0;
    parameter location = "";
    parameter rpath_dynamic = 1'b0;
    parameter rpath_edge = 1'b0;
    parameter rpath_init = 1'b0;
    parameter rpath_load = 1'b0;
    parameter rpath_mode = 4'b0000;
    parameter rpath_sync = 1'b0;
    parameter symbol = "";
    parameter tpath_mode = 2'b00;
    parameter variant = "";
endmodule

(* blackbox *)
module NX_IOM_DRIVER_U(EI1, EI2, EI3, EI4, EI5, EI6, EI7, EI8, EL, ER, CI1, CL, CR, RI, RL, RR, CO, CTI, CTO, EO, RO1
, RO2, RO3, RO4, RO5, RO6, RO7, RO8, LINK);
    input CI1;
    input CL;
    output CO;
    input CR;
    input CTI;
    output CTO;
    input EI1;
    input EI2;
    input EI3;
    input EI4;
    input EI5;
    input EI6;
    input EI7;
    input EI8;
    input EL;
    output EO;
    input ER;
    inout [41:0] LINK;
    input RI;
    input RL;
    output RO1;
    output RO2;
    output RO3;
    output RO4;
    output RO5;
    output RO6;
    output RO7;
    output RO8;
    input RR;
    parameter chained = 1'b0;
    parameter cpath_edge = 1'b0;
    parameter cpath_init = 1'b0;
    parameter cpath_inv = 1'b0;
    parameter cpath_load = 1'b0;
    parameter cpath_mode = 4'b0000;
    parameter cpath_sync = 1'b0;
    parameter cpath_type = 1'b0;
    parameter epath_dynamic = 1'b0;
    parameter epath_edge = 1'b0;
    parameter epath_init = 1'b0;
    parameter epath_load = 1'b0;
    parameter epath_mode = 4'b0000;
    parameter epath_sync = 1'b0;
    parameter epath_type = 1'b0;
    parameter location = "";
    parameter rpath_dynamic = 1'b0;
    parameter rpath_edge = 1'b0;
    parameter rpath_init = 1'b0;
    parameter rpath_load = 1'b0;
    parameter rpath_mode = 4'b0000;
    parameter rpath_sync = 1'b0;
    parameter rpath_type = 1'b0;
    parameter symbol = "";
    parameter tpath_mode = 1'b0;
endmodule

(* blackbox *)
module NX_IOM_SERDES(RTCK, WRCK, WTCK, RRCK, TRST, RRST, CTCK, DCK, DRL, DIG, FZ, FLD, FLG, DS, DRA, DRI, DRO, DID, LINKN, LINKP);
    input CTCK;
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINKN;
    inout [41:0] LINKP;
    input RRCK;
    input RRST;
    input RTCK;
    input TRST;
    input WRCK;
    input WTCK;
    parameter data_size = 5;
    parameter location = "";
endmodule

(* blackbox *)
module NX_IOM_SERDES_M(RTCK, WRCK, WTCK, RRCK, TRST, RRST, CTCK, DCK, DRL, DIG, FZ, FLD, FLG, DS, DRA, DRI, DRO, DID, LINKN, LINKP);
    input CTCK;
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINKN;
    inout [41:0] LINKP;
    input RRCK;
    input RRST;
    input RTCK;
    input TRST;
    input WRCK;
    input WTCK;
    parameter data_size = 5;
    parameter location = "";
endmodule

(* blackbox *)
module NX_IOM_SERDES_U(FCK, SCK, LDRN, DRWDS, DRWEN, DRE, FZ, ALD, ALT, FLD, FLG, LINK, DRA, DRI, DRO, DID, DRIN, DRDN, FA, DRON);
    output ALD;
    output ALT;
    output [5:0] DID;
    input [3:0] DRA;
    input [2:0] DRDN;
    input DRE;
    input [5:0] DRI;
    input [2:0] DRIN;
    output [5:0] DRO;
    input [2:0] DRON;
    input DRWDS;
    input DRWEN;
    input [5:0] FA;
    input FCK;
    output FLD;
    output FLG;
    input FZ;
    input LDRN;
    inout [41:0] LINK;
    input SCK;
    parameter data_size = 5;
    parameter location = "";
endmodule

//(* blackbox *)
//module NX_LUT(I1, I2, I3, I4, O);
//    input I1;
//    input I2;
//    input I3;
//    input I4;
//    output O;
//    parameter lut_table = 16'b0000000000000000;
//endmodule

(* blackbox *)
module NX_RAM(ACK, ACKC, ACKD, ACKR, BCK, BCKC, BCKD, BCKR, AI1, AI2, AI3, AI4, AI5, AI6, AI7, AI8, AI9, AI10, AI11, AI12, AI13
, AI14, AI15, AI16, AI17, AI18, AI19, AI20, AI21, AI22, AI23, AI24, BI1, BI2, BI3, BI4, BI5, BI6, BI7, BI8, BI9, BI10
, BI11, BI12, BI13, BI14, BI15, BI16, BI17, BI18, BI19, BI20, BI21, BI22, BI23, BI24, ACOR, AERR, BCOR, BERR, AO1, AO2, AO3
, AO4, AO5, AO6, AO7, AO8, AO9, AO10, AO11, AO12, AO13, AO14, AO15, AO16, AO17, AO18, AO19, AO20, AO21, AO22, AO23, AO24
, BO1, BO2, BO3, BO4, BO5, BO6, BO7, BO8, BO9, BO10, BO11, BO12, BO13, BO14, BO15, BO16, BO17, BO18, BO19, BO20, BO21
, BO22, BO23, BO24, AA1, AA2, AA3, AA4, AA5, AA6, AA7, AA8, AA9, AA10, AA11, AA12, AA13, AA14, AA15, AA16, ACS, AWE
, AR, BA1, BA2, BA3, BA4, BA5, BA6, BA7, BA8, BA9, BA10, BA11, BA12, BA13, BA14, BA15, BA16, BCS, BWE, BR);
    input AA1;
    input AA10;
    input AA11;
    input AA12;
    input AA13;
    input AA14;
    input AA15;
    input AA16;
    input AA2;
    input AA3;
    input AA4;
    input AA5;
    input AA6;
    input AA7;
    input AA8;
    input AA9;
    input ACK;
    input ACKC;
    input ACKD;
    input ACKR;
    output ACOR;
    input ACS;
    output AERR;
    input AI1;
    input AI10;
    input AI11;
    input AI12;
    input AI13;
    input AI14;
    input AI15;
    input AI16;
    input AI17;
    input AI18;
    input AI19;
    input AI2;
    input AI20;
    input AI21;
    input AI22;
    input AI23;
    input AI24;
    input AI3;
    input AI4;
    input AI5;
    input AI6;
    input AI7;
    input AI8;
    input AI9;
    output AO1;
    output AO10;
    output AO11;
    output AO12;
    output AO13;
    output AO14;
    output AO15;
    output AO16;
    output AO17;
    output AO18;
    output AO19;
    output AO2;
    output AO20;
    output AO21;
    output AO22;
    output AO23;
    output AO24;
    output AO3;
    output AO4;
    output AO5;
    output AO6;
    output AO7;
    output AO8;
    output AO9;
    input AR;
    input AWE;
    input BA1;
    input BA10;
    input BA11;
    input BA12;
    input BA13;
    input BA14;
    input BA15;
    input BA16;
    input BA2;
    input BA3;
    input BA4;
    input BA5;
    input BA6;
    input BA7;
    input BA8;
    input BA9;
    input BCK;
    input BCKC;
    input BCKD;
    input BCKR;
    output BCOR;
    input BCS;
    output BERR;
    input BI1;
    input BI10;
    input BI11;
    input BI12;
    input BI13;
    input BI14;
    input BI15;
    input BI16;
    input BI17;
    input BI18;
    input BI19;
    input BI2;
    input BI20;
    input BI21;
    input BI22;
    input BI23;
    input BI24;
    input BI3;
    input BI4;
    input BI5;
    input BI6;
    input BI7;
    input BI8;
    input BI9;
    output BO1;
    output BO10;
    output BO11;
    output BO12;
    output BO13;
    output BO14;
    output BO15;
    output BO16;
    output BO17;
    output BO18;
    output BO19;
    output BO2;
    output BO20;
    output BO21;
    output BO22;
    output BO23;
    output BO24;
    output BO3;
    output BO4;
    output BO5;
    output BO6;
    output BO7;
    output BO8;
    output BO9;
    input BR;
    input BWE;
    parameter mcka_edge = 1'b0;
    parameter mckb_edge = 1'b0;
    parameter mem_ctxt = "";
    parameter pcka_edge = 1'b0;
    parameter pckb_edge = 1'b0;
    parameter pipe_ia = 1'b0;
    parameter pipe_ib = 1'b0;
    parameter pipe_oa = 1'b0;
    parameter pipe_ob = 1'b0;
    parameter raw_config0 = 4'b0000;
    parameter raw_config1 = 16'b0000000000000000;
    parameter raw_l_enable = 1'b0;
    parameter raw_l_extend = 4'b0000;
    parameter raw_u_enable = 1'b0;
    parameter raw_u_extend = 8'b00000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_RAM_SLOWECC_1K_36_1r1w(ACK, BCK, ACOR, AERR, ACS, AWE, AR, BCS, BWE, BR, AO, AI, AA);
    input [9:0] AA;
    input ACK;
    output ACOR;
    input ACS;
    output AERR;
    input [35:0] AI;
    output [35:0] AO;
    input AR;
    input AWE;
    input BCK;
    input BCS;
    input BR;
    input BWE;
    parameter mem_ctxt = "";
endmodule

(* blackbox *)
module NX_RAM_WRAP(ACK, ACKD, ACKR, BCK, BCKD, BCKR, ACOR, AERR, BCOR, BERR, ACS, AWE, AR, BCS, BWE, BR, BI, AO, BO, AI, AA
, BA);
    input [15:0] AA;
    input ACK;
    input ACKD;
    input ACKR;
    output ACOR;
    input ACS;
    output AERR;
    input [23:0] AI;
    output [23:0] AO;
    input AR;
    input AWE;
    input [15:0] BA;
    input BCK;
    input BCKD;
    input BCKR;
    output BCOR;
    input BCS;
    output BERR;
    input [23:0] BI;
    output [23:0] BO;
    input BR;
    input BWE;
    parameter mcka_edge = 1'b0;
    parameter mckb_edge = 1'b0;
    parameter mem_ctxt = "";
    parameter pcka_edge = 1'b0;
    parameter pckb_edge = 1'b0;
    parameter pipe_ia = 1'b0;
    parameter pipe_ib = 1'b0;
    parameter pipe_oa = 1'b0;
    parameter pipe_ob = 1'b0;
    parameter raw_config0 = 4'b0000;
    parameter raw_config1 = 16'b0000000000000000;
    parameter raw_l_enable = 1'b0;
    parameter raw_l_extend = 4'b0000;
    parameter raw_u_enable = 1'b0;
    parameter raw_u_extend = 8'b00000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_SER(FCK, SCK, R, IO, DCK, DRL, I, DS, DRA, DRI, DRO, DID);
    input DCK;
    output [5:0] DID;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    input FCK;
    input [4:0] I;
    output IO;
    input R;
    input SCK;
    parameter data_size = 5;
    parameter differential = "";
    parameter drive = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter slewRate = "";
    parameter spath_dynamic = 1'b0;
    parameter standard = "";
endmodule

(* blackbox *)
module NX_SERDES(FCK, SCK, RTX, RRX, CI, CCK, CL, CR, IO, DCK, DRL, DIG, FZ, FLD, FLG, I, O, DS, DRA, DRI, DRO
, DID);
    input CCK;
    input CI;
    input CL;
    input CR;
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    input FCK;
    output FLD;
    output FLG;
    input FZ;
    input [4:0] I;
    inout IO;
    output [4:0] O;
    input RRX;
    input RTX;
    input SCK;
    parameter cpath_registered = 1'b0;
    parameter data_size = 5;
    parameter differential = "";
    parameter dpath_dynamic = 1'b0;
    parameter drive = "";
    parameter inputDelayLine = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter slewRate = "";
    parameter spath_dynamic = 1'b0;
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule
