// ---------------------------------------

module \$__ABC_DPR16X4_COMB (input [3:0] A, S, output [3:0] Y);
    assign Y = A;
endmodule
