module test (
    input ia,
    output oa,
    input [0:0] ib,
    output [0:0] ob,
    input [3:0] ic,
    output [3:0] oc
    );

assign oa = ia;
assign ob = ib;
assign oc = ic;

endmodule
