module my_module(
    input a,
    input b,
    output y
);
   // Perform AND
   assign y = a & b;

endmodule
