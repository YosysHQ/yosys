module sub #(parameter d=1) (input in, output out);
    assign out = in;
endmodule
