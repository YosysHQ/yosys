module test(input in, output [1:0] out);
assign out[0] = in;
assign out[1] = in;
endmodule
