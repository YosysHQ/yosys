module unpacked_arrays;
  reg array_range [0:7];
  reg array_size [8];
endmodule
