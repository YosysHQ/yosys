module sub;
    sub _TECHMAP_REPLACE_ ();
    bar f0();
endmodule
