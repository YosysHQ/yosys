(* blackbox *)
module AND(input [7:0] A, B, output [7:0] Y);
endmodule

(* blackbox *)
module ALU(input [7:0] A, B, output [7:0] Y);
parameter MODE = "";
endmodule
