module test(in, out, io, vin, vout, vio);
input in;
output out;
inout io;
input [3:0] vin;
output [3:0] vout;
inout [0:3] vio;
endmodule
