module test(input in, output reg out);

always @(in)
    out = in;
endmodule	
