module C7552_lev2(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, 
	pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, 
	pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, 
	pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, 
	pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, 
	pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, 
	pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, 
	pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, 
	pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, 
	pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, 
	pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, 
	pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, 
	pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, 
	pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, 
	pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, 
	pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, 
	pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, 
	pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, 
	pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, 
	pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, 
	pi200, pi201, pi202, pi203, pi204, pi205, pi206, po000, po001, po002, 
	po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, 
	po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, 
	po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, 
	po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, 
	po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, 
	po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, 
	po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, 
	po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, 
	po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, 
	po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, 
	po103, po104, po105, po106, po107);

input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, 
	pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, 
	pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, 
	pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, 
	pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, 
	pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, 
	pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, 
	pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, 
	pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, 
	pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, 
	pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, 
	pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, 
	pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, 
	pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, 
	pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, 
	pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, 
	pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, 
	pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, 
	pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, 
	pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, 
	pi200, pi201, pi202, pi203, pi204, pi205, pi206;

output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, 
	po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, 
	po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, 
	po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, 
	po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, 
	po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, 
	po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, 
	po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, 
	po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, 
	po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, 
	po100, po101, po102, po103, po104, po105, po106, po107;

wire n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
	n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, 
	n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
	n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, 
	n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
	n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
	n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
	n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
	n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, 
	n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
	n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
	n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, 
	n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, 
	n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
	n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, 
	n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
	n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
	n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
	n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, 
	n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
	n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, 
	n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, 
	n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, 
	n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, 
	n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, 
	n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
	n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
	n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
	n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
	n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
	n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
	n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
	n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
	n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
	n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
	n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
	n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
	n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
	n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
	n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
	n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
	n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
	n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, 
	n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, 
	n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
	n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
	n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
	n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, 
	n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
	n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
	n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
	n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
	n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
	n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
	n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, 
	n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
	n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
	n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
	n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
	n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
	n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
	n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
	n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
	n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
	n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
	n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
	n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, 
	n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
	n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, 
	n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
	n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
	n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
	n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
	n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, 
	n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, 
	n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
	n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, 
	n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, 
	n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, 
	n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, 
	n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, 
	n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
	n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, 
	n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, 
	n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, 
	n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
	n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
	n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
	n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
	n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
	n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
	n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
	n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
	n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
	n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
	n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
	n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
	n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
	n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
	n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
	n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
	n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, 
	n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
	n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, 
	n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, 
	n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
	n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
	n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
	n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
	n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, 
	n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, 
	n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, 
	n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
	n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, 
	n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, 
	n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, 
	n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, 
	n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, 
	n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, 
	n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, 
	n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, 
	n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, 
	n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, 
	n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, 
	n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, 
	n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, 
	n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, 
	n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, 
	n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, 
	n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, 
	n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, 
	n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, 
	n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, 
	n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, 
	n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, 
	n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, 
	n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, 
	n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, 
	n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, 
	n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, 
	n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, 
	n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, 
	n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, 
	n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, 
	n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, 
	n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, 
	n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, 
	n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, 
	n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, 
	n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, 
	n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, 
	n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
	n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, 
	n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, 
	n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, 
	n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, 
	n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, 
	n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, 
	n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, 
	n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, 
	n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, 
	n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, 
	n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, 
	n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, 
	n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, 
	n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, 
	n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, 
	n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, 
	n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, 
	n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, 
	n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, 
	n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, 
	n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, 
	n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, 
	n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, 
	n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, 
	n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, 
	n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, 
	n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, 
	n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, 
	n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, 
	n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, 
	n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, 
	n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, 
	n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, 
	n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, 
	n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, 
	n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, 
	n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, 
	n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, 
	n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, 
	n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, 
	n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, 
	n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, 
	n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, 
	n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, 
	n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, 
	n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, 
	n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, 
	n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, 
	n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, 
	n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, 
	n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, 
	n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, 
	n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, 
	n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, 
	n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, 
	n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, 
	n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, 
	n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, 
	n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, 
	n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, 
	n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, 
	n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, 
	n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, 
	n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, 
	n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, 
	n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, 
	n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, 
	n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, 
	n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, 
	n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, 
	n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, 
	n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, 
	n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, 
	n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, 
	n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, 
	n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, 
	n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, 
	n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, 
	n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, 
	n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, 
	n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, 
	n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, 
	n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, 
	n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, 
	n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, 
	n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, 
	n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, 
	n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, 
	n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, 
	n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, 
	n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, 
	n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, 
	n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, 
	n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, 
	n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, 
	n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, 
	n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, 
	n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, 
	n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, 
	n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, 
	n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, 
	n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, 
	n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, 
	n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, 
	n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, 
	n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, 
	n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, 
	n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, 
	n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, 
	n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, 
	n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, 
	n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, 
	n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
	n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, 
	n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, 
	n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, 
	n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, 
	n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
	n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, 
	n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, 
	n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, 
	n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, 
	n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, 
	n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
	n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
	n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
	n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
	n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
	n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
	n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, 
	n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, 
	n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
	n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, 
	n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
	n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, 
	n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
	n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
	n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, 
	n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, 
	n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
	n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, 
	n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
	n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, 
	n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
	n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, 
	n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, 
	n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
	n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
	n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, 
	n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, 
	n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, 
	n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
	n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, 
	n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, 
	n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, 
	n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, 
	n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
	n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, 
	n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, 
	n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, 
	n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, 
	n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
	n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, 
	n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
	n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
	n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
	n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
	n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
	n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, 
	n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, 
	n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, 
	n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
	n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
	n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
	n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, 
	n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
	n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
	n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, 
	n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
	n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
	n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
	n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
	n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, 
	n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
	n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
	n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
	n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
	n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
	n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
	n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
	n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
	n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
	n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
	n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
	n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
	n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
	n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
	n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
	n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
	n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
	n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
	n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
	n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
	n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
	n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
	n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
	n6402, n6403, n6404, n6405;

assign po001 = pi187;

assign po015 = po003;

assign po004 = pi106;

assign po009 = pi136;

assign po010 = pi022;

assign po011 = pi112;

assign po005 = po012;

assign po013 = pi062;

assign po014 = pi123;

assign po101 = po023;

assign po067 = po023;

assign po066 = po023;

assign po023 = pi119;

assign po024 = pi152;

assign po025 = pi125;

assign po027 = pi102;

assign po028 = pi031;

assign po031 = pi155;

assign po065 = po034;

assign po035 = pi182;

assign po036 = pi023;

assign po038 = pi071;

assign po039 = pi015;

assign po040 = pi132;

assign po044 = pi044;

assign po052 = pi048;

assign po057 = pi117;

assign po059 = pi091;

assign po063 = pi000;

assign po064 = pi194;

assign po069 = pi147;

assign po070 = pi002;

assign po071 = pi080;

assign po072 = pi188;

assign po018 = po074;

assign po021 = po074;

assign po079 = pi084;

assign po082 = pi144;

assign po084 = pi199;

assign po085 = pi066;

assign po091 = pi008;

assign po092 = pi154;

assign po099 = pi042;

assign po102 = pi179;

assign po103 = pi145;

assign po104 = pi127;

assign po106 = pi105;

assign po107 = pi029;

assign po020 = po041;

assign po032 = po007;

assign po089 = po076;

assign po054 = po076;

  OR2 U2865 ( .A(n2822), .B(n2823), .Z(po100));
  AN2 U2866 ( .A(n2824), .B(pi192), .Z(n2823));
  OR2 U2867 ( .A(n2825), .B(n2826), .Z(n2824));
  AN2 U2868 ( .A(n2827), .B(n2828), .Z(n2826));
  IV2 U2869 ( .A(n2829), .Z(n2825));
  OR2 U2870 ( .A(n2828), .B(n2827), .Z(n2829));
  OR2 U2871 ( .A(n2830), .B(n2831), .Z(n2827));
  AN2 U2872 ( .A(n2832), .B(n2833), .Z(n2831));
  AN2 U2873 ( .A(n2834), .B(n2835), .Z(n2830));
  AN2 U2874 ( .A(n2836), .B(n2837), .Z(n2822));
  OR2 U2875 ( .A(n2838), .B(n2839), .Z(n2836));
  AN2 U2876 ( .A(n2840), .B(n2828), .Z(n2839));
  IV2 U2877 ( .A(n2841), .Z(n2838));
  OR2 U2878 ( .A(n2828), .B(n2840), .Z(n2841));
  OR2 U2879 ( .A(n2842), .B(n2843), .Z(n2840));
  AN2 U2880 ( .A(n2844), .B(n2845), .Z(n2843));
  AN2 U2881 ( .A(n2846), .B(n2847), .Z(n2842));
  AN2 U2882 ( .A(n2848), .B(n2849), .Z(n2828));
  IV2 U2883 ( .A(n2850), .Z(n2849));
  AN2 U2884 ( .A(n2851), .B(n2852), .Z(n2850));
  OR2 U2885 ( .A(n2852), .B(n2851), .Z(n2848));
  OR2 U2886 ( .A(n2853), .B(n2854), .Z(n2851));
  AN2 U2887 ( .A(n2855), .B(n2856), .Z(n2854));
  IV2 U2888 ( .A(n2857), .Z(n2853));
  OR2 U2889 ( .A(n2856), .B(n2855), .Z(n2857));
  IV2 U2890 ( .A(n2858), .Z(n2855));
  OR2 U2891 ( .A(n2859), .B(n2860), .Z(n2858));
  AN2 U2892 ( .A(n2861), .B(n2862), .Z(n2859));
  OR2 U2893 ( .A(n2863), .B(n2864), .Z(n2856));
  OR2 U2894 ( .A(n2865), .B(n2866), .Z(n2864));
  AN2 U2895 ( .A(pi192), .B(n2867), .Z(n2866));
  OR2 U2896 ( .A(n2868), .B(n2869), .Z(n2867));
  OR2 U2897 ( .A(n2870), .B(n2871), .Z(n2869));
  AN2 U2898 ( .A(n2872), .B(n2873), .Z(n2871));
  AN2 U2899 ( .A(n2862), .B(n2874), .Z(n2872));
  OR2 U2900 ( .A(n2875), .B(n2876), .Z(n2874));
  AN2 U2901 ( .A(n2877), .B(n2878), .Z(n2875));
  AN2 U2902 ( .A(n2879), .B(n2880), .Z(n2870));
  AN2 U2903 ( .A(n2881), .B(n2882), .Z(n2868));
  OR2 U2904 ( .A(n2883), .B(n2884), .Z(n2881));
  AN2 U2905 ( .A(n2885), .B(n2886), .Z(n2884));
  AN2 U2906 ( .A(n2879), .B(n2887), .Z(n2883));
  IV2 U2907 ( .A(n2873), .Z(n2879));
  OR2 U2908 ( .A(n2888), .B(n2889), .Z(n2873));
  AN2 U2909 ( .A(n2890), .B(n2891), .Z(n2889));
  AN2 U2910 ( .A(n2892), .B(n2886), .Z(n2888));
  AN2 U2911 ( .A(n2893), .B(n2837), .Z(n2865));
  OR2 U2912 ( .A(n2894), .B(n2895), .Z(n2893));
  OR2 U2913 ( .A(n2896), .B(n2897), .Z(n2895));
  OR2 U2914 ( .A(n2898), .B(n2899), .Z(n2897));
  AN2 U2915 ( .A(n2900), .B(n2901), .Z(n2899));
  AN2 U2916 ( .A(n2902), .B(n2903), .Z(n2900));
  OR2 U2917 ( .A(n2904), .B(n2905), .Z(n2903));
  OR2 U2918 ( .A(n2906), .B(n2907), .Z(n2905));
  AN2 U2919 ( .A(n2890), .B(n2908), .Z(n2907));
  AN2 U2920 ( .A(n2909), .B(n2886), .Z(n2906));
  AN2 U2921 ( .A(n2910), .B(pi082), .Z(n2909));
  AN2 U2922 ( .A(pi200), .B(n2911), .Z(n2898));
  OR2 U2923 ( .A(n2912), .B(n2913), .Z(n2911));
  OR2 U2924 ( .A(n2914), .B(n2915), .Z(n2913));
  AN2 U2925 ( .A(n2916), .B(n2890), .Z(n2915));
  AN2 U2926 ( .A(n2910), .B(n2917), .Z(n2916));
  OR2 U2927 ( .A(n2918), .B(n2919), .Z(n2917));
  AN2 U2928 ( .A(n2920), .B(n2886), .Z(n2914));
  OR2 U2929 ( .A(n2921), .B(n2922), .Z(n2920));
  OR2 U2930 ( .A(n2923), .B(n2924), .Z(n2922));
  AN2 U2931 ( .A(n2918), .B(n2860), .Z(n2924));
  AN2 U2932 ( .A(n2925), .B(n2926), .Z(n2923));
  OR2 U2933 ( .A(n2927), .B(n2928), .Z(n2926));
  AN2 U2934 ( .A(n2844), .B(n2929), .Z(n2928));
  AN2 U2935 ( .A(n2930), .B(n2931), .Z(n2927));
  OR2 U2936 ( .A(n2932), .B(n2933), .Z(n2921));
  AN2 U2937 ( .A(n2934), .B(n2935), .Z(n2933));
  AN2 U2938 ( .A(n2936), .B(n2910), .Z(n2934));
  AN2 U2939 ( .A(n2937), .B(n2938), .Z(n2932));
  AN2 U2940 ( .A(n2929), .B(n2939), .Z(n2937));
  AN2 U2941 ( .A(n2935), .B(n2940), .Z(n2912));
  OR2 U2942 ( .A(n2904), .B(n2941), .Z(n2940));
  AN2 U2943 ( .A(n2890), .B(n2942), .Z(n2941));
  AN2 U2944 ( .A(n2943), .B(n2944), .Z(n2942));
  OR2 U2945 ( .A(n2945), .B(n2946), .Z(n2944));
  IV2 U2946 ( .A(n2910), .Z(n2945));
  OR2 U2947 ( .A(n2936), .B(n2947), .Z(n2943));
  IV2 U2948 ( .A(n2948), .Z(n2904));
  OR2 U2949 ( .A(n2949), .B(n2939), .Z(n2948));
  AN2 U2950 ( .A(n2950), .B(n2951), .Z(n2949));
  OR2 U2951 ( .A(n2890), .B(n2947), .Z(n2951));
  OR2 U2952 ( .A(n2929), .B(n2886), .Z(n2950));
  AN2 U2953 ( .A(n2952), .B(n2953), .Z(n2896));
  AN2 U2954 ( .A(n2954), .B(n2955), .Z(n2953));
  OR2 U2955 ( .A(n2956), .B(n2957), .Z(n2955));
  AN2 U2956 ( .A(n2890), .B(n2958), .Z(n2956));
  OR2 U2957 ( .A(n2959), .B(n2960), .Z(n2958));
  OR2 U2958 ( .A(pi082), .B(n2961), .Z(n2954));
  AN2 U2959 ( .A(n2901), .B(n2886), .Z(n2961));
  AN2 U2960 ( .A(n2910), .B(n2962), .Z(n2952));
  AN2 U2961 ( .A(n2947), .B(n2862), .Z(n2910));
  OR2 U2962 ( .A(n2963), .B(n2964), .Z(n2894));
  AN2 U2963 ( .A(n2965), .B(n2890), .Z(n2964));
  AN2 U2964 ( .A(n2929), .B(n2966), .Z(n2965));
  OR2 U2965 ( .A(n2967), .B(n2968), .Z(n2966));
  AN2 U2966 ( .A(n2969), .B(n2901), .Z(n2967));
  OR2 U2967 ( .A(n2970), .B(n2971), .Z(n2969));
  OR2 U2968 ( .A(n2972), .B(n2973), .Z(n2971));
  AN2 U2969 ( .A(n2902), .B(n2962), .Z(n2973));
  AN2 U2970 ( .A(n2974), .B(n2957), .Z(n2972));
  AN2 U2971 ( .A(pi082), .B(po031), .Z(n2970));
  AN2 U2972 ( .A(n2975), .B(n2886), .Z(n2963));
  OR2 U2973 ( .A(n2976), .B(n2977), .Z(n2975));
  AN2 U2974 ( .A(n2968), .B(n2947), .Z(n2977));
  AN2 U2975 ( .A(n2978), .B(n2979), .Z(n2968));
  OR2 U2976 ( .A(n2980), .B(n2981), .Z(n2979));
  AN2 U2977 ( .A(n2982), .B(n2931), .Z(n2980));
  AN2 U2978 ( .A(n2983), .B(n2929), .Z(n2976));
  AN2 U2979 ( .A(n2984), .B(n2936), .Z(n2983));
  AN2 U2980 ( .A(n2974), .B(n2901), .Z(n2984));
  OR2 U2981 ( .A(n2985), .B(n2986), .Z(n2863));
  AN2 U2982 ( .A(n2987), .B(n2890), .Z(n2986));
  AN2 U2983 ( .A(n2988), .B(n2989), .Z(n2987));
  AN2 U2984 ( .A(n2990), .B(n2962), .Z(n2989));
  AN2 U2985 ( .A(n2862), .B(n2877), .Z(n2988));
  AN2 U2986 ( .A(n2991), .B(n2886), .Z(n2985));
  OR2 U2987 ( .A(n2992), .B(n2993), .Z(n2991));
  AN2 U2988 ( .A(n2994), .B(n2995), .Z(n2993));
  AN2 U2989 ( .A(n2990), .B(n2901), .Z(n2995));
  AN2 U2990 ( .A(n2996), .B(n2974), .Z(n2994));
  OR2 U2991 ( .A(po031), .B(n2930), .Z(n2996));
  AN2 U2992 ( .A(n2997), .B(n2860), .Z(n2992));
  AN2 U2993 ( .A(n2998), .B(n2930), .Z(n2860));
  AN2 U2994 ( .A(n2877), .B(n2999), .Z(n2997));
  IV2 U2995 ( .A(n2882), .Z(n2877));
  AN2 U2996 ( .A(n3000), .B(n3001), .Z(n2852));
  OR2 U2997 ( .A(n3002), .B(n2925), .Z(n3001));
  OR2 U2998 ( .A(n3003), .B(n3004), .Z(n3000));
  IV2 U2999 ( .A(n3002), .Z(n3004));
  OR2 U3000 ( .A(n3005), .B(n3006), .Z(n3002));
  AN2 U3001 ( .A(n3007), .B(n3008), .Z(n3006));
  OR2 U3002 ( .A(n3009), .B(n3010), .Z(n3008));
  AN2 U3003 ( .A(n3011), .B(n3012), .Z(n3009));
  AN2 U3004 ( .A(n3013), .B(n3014), .Z(n3007));
  OR2 U3005 ( .A(n3015), .B(n3016), .Z(n3014));
  IV2 U3006 ( .A(n3017), .Z(n3016));
  OR2 U3007 ( .A(n3017), .B(n3018), .Z(n3013));
  OR2 U3008 ( .A(n3019), .B(n3020), .Z(n3017));
  AN2 U3009 ( .A(n3021), .B(n3022), .Z(n3020));
  OR2 U3010 ( .A(n3023), .B(n3024), .Z(n3022));
  OR2 U3011 ( .A(n3025), .B(n3026), .Z(n3024));
  OR2 U3012 ( .A(n3027), .B(n3028), .Z(n3026));
  AN2 U3013 ( .A(po010), .B(n3029), .Z(n3028));
  AN2 U3014 ( .A(n3030), .B(pi192), .Z(n3027));
  AN2 U3015 ( .A(n3031), .B(n3032), .Z(n3030));
  OR2 U3016 ( .A(n3033), .B(n3034), .Z(n3032));
  AN2 U3017 ( .A(n3035), .B(n3036), .Z(n3034));
  AN2 U3018 ( .A(n3015), .B(n3037), .Z(n3035));
  OR2 U3019 ( .A(n3038), .B(n3039), .Z(n3031));
  OR2 U3020 ( .A(n3040), .B(n3041), .Z(n3039));
  AN2 U3021 ( .A(po010), .B(n3042), .Z(n3040));
  OR2 U3022 ( .A(n3043), .B(n3044), .Z(n3025));
  AN2 U3023 ( .A(n3015), .B(n3045), .Z(n3044));
  OR2 U3024 ( .A(n3046), .B(n3047), .Z(n3045));
  AN2 U3025 ( .A(n3048), .B(n3049), .Z(n3047));
  OR2 U3026 ( .A(n3050), .B(n3051), .Z(n3048));
  AN2 U3027 ( .A(n3052), .B(po070), .Z(n3051));
  AN2 U3028 ( .A(n3053), .B(po099), .Z(n3050));
  AN2 U3029 ( .A(n3054), .B(n3055), .Z(n3046));
  AN2 U3030 ( .A(n3018), .B(n3056), .Z(n3043));
  OR2 U3031 ( .A(n3057), .B(n3058), .Z(n3056));
  OR2 U3032 ( .A(n3059), .B(n3060), .Z(n3058));
  AN2 U3033 ( .A(n3061), .B(n3042), .Z(n3060));
  AN2 U3034 ( .A(n3062), .B(n3063), .Z(n3059));
  AN2 U3035 ( .A(n3064), .B(n3049), .Z(n3062));
  AN2 U3036 ( .A(n3065), .B(n3066), .Z(n3057));
  OR2 U3037 ( .A(n3067), .B(n3068), .Z(n3023));
  OR2 U3038 ( .A(n3069), .B(n3070), .Z(n3068));
  AN2 U3039 ( .A(n3071), .B(n3072), .Z(n3070));
  AN2 U3040 ( .A(n3053), .B(n3073), .Z(n3069));
  OR2 U3041 ( .A(n3074), .B(n3075), .Z(n3067));
  AN2 U3042 ( .A(n3076), .B(n3077), .Z(n3075));
  OR2 U3043 ( .A(n3078), .B(n3079), .Z(n3077));
  AN2 U3044 ( .A(n3080), .B(n3066), .Z(n3078));
  AN2 U3045 ( .A(n3081), .B(n3061), .Z(n3074));
  AN2 U3046 ( .A(n3082), .B(n3038), .Z(n3081));
  AN2 U3047 ( .A(n3083), .B(n3084), .Z(n3019));
  OR2 U3048 ( .A(n3085), .B(n3086), .Z(n3084));
  OR2 U3049 ( .A(n3087), .B(n3088), .Z(n3086));
  OR2 U3050 ( .A(n3089), .B(n3090), .Z(n3088));
  AN2 U3051 ( .A(n3091), .B(n3049), .Z(n3089));
  OR2 U3052 ( .A(n3092), .B(n3093), .Z(n3087));
  AN2 U3053 ( .A(n3015), .B(n3094), .Z(n3093));
  OR2 U3054 ( .A(n3095), .B(n3096), .Z(n3094));
  OR2 U3055 ( .A(n3097), .B(n3098), .Z(n3096));
  AN2 U3056 ( .A(n3099), .B(n3100), .Z(n3098));
  AN2 U3057 ( .A(po010), .B(po070), .Z(n3099));
  AN2 U3058 ( .A(n3101), .B(pi192), .Z(n3097));
  AN2 U3059 ( .A(n3041), .B(n3038), .Z(n3101));
  OR2 U3060 ( .A(n3102), .B(n3103), .Z(n3041));
  AN2 U3061 ( .A(n3104), .B(pi166), .Z(n3103));
  AN2 U3062 ( .A(n3037), .B(n3049), .Z(n3104));
  AN2 U3063 ( .A(n3105), .B(n3106), .Z(n3102));
  OR2 U3064 ( .A(n3107), .B(n3042), .Z(n3105));
  AN2 U3065 ( .A(po010), .B(n3108), .Z(n3107));
  AN2 U3066 ( .A(n3079), .B(n3109), .Z(n3095));
  OR2 U3067 ( .A(n3110), .B(n3111), .Z(n3079));
  AN2 U3068 ( .A(n3071), .B(n3112), .Z(n3111));
  AN2 U3069 ( .A(n3065), .B(n3113), .Z(n3110));
  OR2 U3070 ( .A(n3114), .B(n3066), .Z(n3113));
  AN2 U3071 ( .A(po010), .B(n3115), .Z(n3114));
  AN2 U3072 ( .A(n3018), .B(n3116), .Z(n3092));
  OR2 U3073 ( .A(n3117), .B(n3118), .Z(n3116));
  AN2 U3074 ( .A(n3065), .B(n3119), .Z(n3118));
  AN2 U3075 ( .A(n3063), .B(n3120), .Z(n3117));
  OR2 U3076 ( .A(n3121), .B(n3122), .Z(n3085));
  OR2 U3077 ( .A(n3123), .B(n3124), .Z(n3122));
  AN2 U3078 ( .A(n3125), .B(n3055), .Z(n3124));
  AN2 U3079 ( .A(n3076), .B(n3112), .Z(n3125));
  AN2 U3080 ( .A(n3126), .B(n3127), .Z(n3123));
  AN2 U3081 ( .A(n3033), .B(n3037), .Z(n3126));
  AN2 U3082 ( .A(n3080), .B(n3072), .Z(n3121));
  AN2 U3083 ( .A(n3119), .B(n3018), .Z(n3072));
  AN2 U3084 ( .A(n3128), .B(n3129), .Z(n3005));
  OR2 U3085 ( .A(n3130), .B(n3131), .Z(n3129));
  OR2 U3086 ( .A(n3132), .B(n3133), .Z(n3131));
  AN2 U3087 ( .A(n3134), .B(pi192), .Z(n3133));
  AN2 U3088 ( .A(n3135), .B(n3136), .Z(n3134));
  OR2 U3089 ( .A(n3137), .B(po044), .Z(n3135));
  AN2 U3090 ( .A(n3138), .B(n2886), .Z(n3137));
  AN2 U3091 ( .A(n3139), .B(n2837), .Z(n3132));
  AN2 U3092 ( .A(n3140), .B(n3141), .Z(n3139));
  OR2 U3093 ( .A(n3142), .B(po044), .Z(n3140));
  AN2 U3094 ( .A(n3143), .B(n2886), .Z(n3142));
  AN2 U3095 ( .A(n3144), .B(n3145), .Z(n3130));
  OR2 U3096 ( .A(n3146), .B(n3147), .Z(n3145));
  IV2 U3097 ( .A(n3012), .Z(n3144));
  AN2 U3098 ( .A(n3148), .B(n3149), .Z(n3128));
  OR2 U3099 ( .A(n3150), .B(n3018), .Z(n3149));
  OR2 U3100 ( .A(n3015), .B(n3151), .Z(n3148));
  IV2 U3101 ( .A(n3150), .Z(n3151));
  OR2 U3102 ( .A(n3152), .B(n3153), .Z(n3150));
  AN2 U3103 ( .A(n3021), .B(n3154), .Z(n3153));
  AN2 U3104 ( .A(n3155), .B(n3083), .Z(n3152));
  IV2 U3105 ( .A(n3154), .Z(n3155));
  OR2 U3106 ( .A(n3156), .B(n3157), .Z(n3154));
  OR2 U3107 ( .A(n3091), .B(n3158), .Z(n3157));
  OR2 U3108 ( .A(n3159), .B(n3160), .Z(n3158));
  AN2 U3109 ( .A(n3161), .B(n3049), .Z(n3160));
  OR2 U3110 ( .A(n3162), .B(n3029), .Z(n3161));
  OR2 U3111 ( .A(n3163), .B(n3164), .Z(n3029));
  AN2 U3112 ( .A(po099), .B(n3165), .Z(n3164));
  OR2 U3113 ( .A(n3166), .B(n3167), .Z(n3165));
  OR2 U3114 ( .A(n3168), .B(n3169), .Z(n3167));
  AN2 U3115 ( .A(n3170), .B(pi192), .Z(n3169));
  AN2 U3116 ( .A(n3038), .B(n3171), .Z(n3170));
  AN2 U3117 ( .A(n3054), .B(n2837), .Z(n3168));
  AN2 U3118 ( .A(n3172), .B(n3173), .Z(n3166));
  AN2 U3119 ( .A(n3015), .B(n3109), .Z(n3172));
  AN2 U3120 ( .A(n3100), .B(n3018), .Z(n3163));
  AN2 U3121 ( .A(n3015), .B(n3174), .Z(n3162));
  OR2 U3122 ( .A(n3175), .B(n3176), .Z(n3174));
  AN2 U3123 ( .A(n3054), .B(n3173), .Z(n3176));
  AN2 U3124 ( .A(n3177), .B(n3109), .Z(n3054));
  AN2 U3125 ( .A(n3178), .B(n3064), .Z(n3175));
  AN2 U3126 ( .A(n3038), .B(n3037), .Z(n3178));
  AN2 U3127 ( .A(po010), .B(n3179), .Z(n3159));
  OR2 U3128 ( .A(n3090), .B(n3180), .Z(n3179));
  OR2 U3129 ( .A(n3181), .B(n3182), .Z(n3180));
  AN2 U3130 ( .A(n3053), .B(n3183), .Z(n3182));
  OR2 U3131 ( .A(n3184), .B(n3119), .Z(n3183));
  AN2 U3132 ( .A(pi141), .B(n3015), .Z(n3184));
  AN2 U3133 ( .A(n3109), .B(n3065), .Z(n3053));
  AN2 U3134 ( .A(n3185), .B(n3061), .Z(n3181));
  AN2 U3135 ( .A(n3186), .B(n3038), .Z(n3185));
  OR2 U3136 ( .A(n3187), .B(n3063), .Z(n3186));
  AN2 U3137 ( .A(pi033), .B(n3015), .Z(n3187));
  OR2 U3138 ( .A(n3188), .B(n3189), .Z(n3090));
  AN2 U3139 ( .A(n3190), .B(n3065), .Z(n3189));
  AN2 U3140 ( .A(n3073), .B(n3076), .Z(n3190));
  AN2 U3141 ( .A(n3191), .B(n3061), .Z(n3188));
  AN2 U3142 ( .A(n3082), .B(n3033), .Z(n3191));
  OR2 U3143 ( .A(n3192), .B(n3193), .Z(n3091));
  OR2 U3144 ( .A(n3194), .B(n3195), .Z(n3193));
  AN2 U3145 ( .A(n3052), .B(n3018), .Z(n3195));
  AN2 U3146 ( .A(n3064), .B(n3196), .Z(n3194));
  OR2 U3147 ( .A(n3197), .B(n3198), .Z(n3196));
  AN2 U3148 ( .A(n3082), .B(n3199), .Z(n3198));
  AN2 U3149 ( .A(n3042), .B(n3033), .Z(n3197));
  OR2 U3150 ( .A(n3200), .B(n3201), .Z(n3192));
  AN2 U3151 ( .A(n3173), .B(n3202), .Z(n3201));
  OR2 U3152 ( .A(n3203), .B(n3204), .Z(n3202));
  AN2 U3153 ( .A(n3073), .B(n3205), .Z(n3204));
  AN2 U3154 ( .A(n3076), .B(n3066), .Z(n3203));
  AN2 U3155 ( .A(n3206), .B(po099), .Z(n3200));
  AN2 U3156 ( .A(po070), .B(n3207), .Z(n3206));
  OR2 U3157 ( .A(n3208), .B(n3209), .Z(n3156));
  AN2 U3158 ( .A(n3210), .B(n3055), .Z(n3209));
  AN2 U3159 ( .A(n3076), .B(n3115), .Z(n3210));
  AN2 U3160 ( .A(n3211), .B(n3127), .Z(n3208));
  AN2 U3161 ( .A(n3033), .B(n3108), .Z(n3211));
  OR2 U3162 ( .A(n3212), .B(n3213), .Z(po098));
  AN2 U3163 ( .A(n3214), .B(pi192), .Z(n3213));
  OR2 U3164 ( .A(n3215), .B(n3216), .Z(n3214));
  AN2 U3165 ( .A(n2832), .B(n2901), .Z(n3216));
  IV2 U3166 ( .A(n2835), .Z(n2832));
  AN2 U3167 ( .A(pi200), .B(n2835), .Z(n3215));
  OR2 U3168 ( .A(n2880), .B(n2876), .Z(n2835));
  AN2 U3169 ( .A(n3217), .B(n2837), .Z(n3212));
  OR2 U3170 ( .A(n3218), .B(n3219), .Z(n3217));
  AN2 U3171 ( .A(n3220), .B(n2847), .Z(n3219));
  OR2 U3172 ( .A(n3221), .B(n2902), .Z(n3220));
  AN2 U3173 ( .A(pi200), .B(n2938), .Z(n3221));
  AN2 U3174 ( .A(n2844), .B(n3222), .Z(n3218));
  IV2 U3175 ( .A(n2847), .Z(n2844));
  OR2 U3176 ( .A(n2936), .B(n2978), .Z(n2847));
  OR2 U3177 ( .A(n3223), .B(n3224), .Z(po097));
  AN2 U3178 ( .A(n3225), .B(n3226), .Z(n3224));
  OR2 U3179 ( .A(n3227), .B(n3228), .Z(n3226));
  OR2 U3180 ( .A(n3229), .B(n3230), .Z(n3228));
  OR2 U3181 ( .A(n3231), .B(n3232), .Z(n3230));
  AN2 U3182 ( .A(n3233), .B(n3234), .Z(n3232));
  AN2 U3183 ( .A(n3235), .B(n3236), .Z(n3231));
  OR2 U3184 ( .A(n3237), .B(n3238), .Z(n3227));
  OR2 U3185 ( .A(n3239), .B(n3240), .Z(n3238));
  AN2 U3186 ( .A(n3241), .B(n3242), .Z(n3240));
  AN2 U3187 ( .A(n3243), .B(n3244), .Z(n3239));
  AN2 U3188 ( .A(po082), .B(n3245), .Z(n3237));
  AN2 U3189 ( .A(n3246), .B(n3247), .Z(n3223));
  OR2 U3190 ( .A(n3248), .B(n3249), .Z(n3246));
  AN2 U3191 ( .A(n3250), .B(n3251), .Z(n3249));
  OR2 U3192 ( .A(n3252), .B(n3253), .Z(po096));
  AN2 U3193 ( .A(n3254), .B(n3255), .Z(n3252));
  OR2 U3194 ( .A(n3256), .B(n3257), .Z(n3254));
  AN2 U3195 ( .A(n3258), .B(n3259), .Z(n3256));
  AN2 U3196 ( .A(n3260), .B(n3261), .Z(n3258));
  OR2 U3197 ( .A(n3262), .B(n3263), .Z(n3260));
  AN2 U3198 ( .A(n3264), .B(n3265), .Z(n3262));
  OR2 U3199 ( .A(n3266), .B(n3267), .Z(po095));
  OR2 U3200 ( .A(n3268), .B(n3269), .Z(n3267));
  AN2 U3201 ( .A(n3270), .B(n3119), .Z(n3269));
  OR2 U3202 ( .A(n3271), .B(n3272), .Z(n3270));
  AN2 U3203 ( .A(n3273), .B(n2837), .Z(n3272));
  AN2 U3204 ( .A(n3065), .B(n3274), .Z(n3271));
  AN2 U3205 ( .A(n3063), .B(n3275), .Z(n3268));
  OR2 U3206 ( .A(n3276), .B(n3277), .Z(n3275));
  AN2 U3207 ( .A(n3273), .B(pi192), .Z(n3277));
  AN2 U3208 ( .A(n3061), .B(n3274), .Z(n3276));
  OR2 U3209 ( .A(n3278), .B(n3279), .Z(n3266));
  AN2 U3210 ( .A(n3280), .B(n3281), .Z(n3279));
  OR2 U3211 ( .A(n3282), .B(n3100), .Z(n3281));
  AN2 U3212 ( .A(n3283), .B(n3284), .Z(n3278));
  OR2 U3213 ( .A(n3285), .B(n3052), .Z(n3283));
  AN2 U3214 ( .A(n3286), .B(n3287), .Z(n3052));
  AN2 U3215 ( .A(po099), .B(n3207), .Z(n3285));
  AN2 U3216 ( .A(n3288), .B(n3289), .Z(po094));
  OR2 U3217 ( .A(n3290), .B(n3291), .Z(n3289));
  OR2 U3218 ( .A(n3234), .B(n3292), .Z(n3288));
  OR2 U3219 ( .A(n3293), .B(n3294), .Z(po093));
  AN2 U3220 ( .A(n3295), .B(n3296), .Z(n3294));
  OR2 U3221 ( .A(n3297), .B(n3298), .Z(n3296));
  AN2 U3222 ( .A(n3299), .B(n3300), .Z(n3297));
  AN2 U3223 ( .A(n3301), .B(n3302), .Z(n3293));
  IV2 U3224 ( .A(n3303), .Z(n3302));
  AN2 U3225 ( .A(n3304), .B(n3299), .Z(n3303));
  OR2 U3226 ( .A(n3305), .B(n3306), .Z(n3299));
  OR2 U3227 ( .A(n3300), .B(n3298), .Z(n3304));
  AN2 U3228 ( .A(n3305), .B(n3306), .Z(n3298));
  OR2 U3229 ( .A(n3307), .B(n3308), .Z(po090));
  OR2 U3230 ( .A(n3309), .B(n3310), .Z(n3308));
  AN2 U3231 ( .A(n3311), .B(n3312), .Z(n3310));
  AN2 U3232 ( .A(n3313), .B(n3314), .Z(n3309));
  OR2 U3233 ( .A(n3315), .B(n3316), .Z(n3313));
  OR2 U3234 ( .A(n3317), .B(n3318), .Z(n3316));
  AN2 U3235 ( .A(n3319), .B(n3320), .Z(n3315));
  OR2 U3236 ( .A(n3321), .B(n3322), .Z(n3319));
  OR2 U3237 ( .A(n3323), .B(n3324), .Z(n3307));
  AN2 U3238 ( .A(n3325), .B(n3326), .Z(n3324));
  AN2 U3239 ( .A(n3327), .B(n3328), .Z(n3323));
  OR2 U3240 ( .A(n3329), .B(n3330), .Z(n3327));
  OR2 U3241 ( .A(n3331), .B(n3332), .Z(po088));
  IV2 U3242 ( .A(n3333), .Z(n3332));
  OR2 U3243 ( .A(n3334), .B(n3335), .Z(n3333));
  AN2 U3244 ( .A(n3335), .B(n3334), .Z(n3331));
  AN2 U3245 ( .A(n3336), .B(n3337), .Z(n3334));
  OR2 U3246 ( .A(n3338), .B(n3339), .Z(n3337));
  IV2 U3247 ( .A(n3340), .Z(n3338));
  OR2 U3248 ( .A(n3341), .B(n3340), .Z(n3336));
  OR2 U3249 ( .A(n3342), .B(n3343), .Z(n3340));
  AN2 U3250 ( .A(n3291), .B(n3250), .Z(n3343));
  AN2 U3251 ( .A(n3344), .B(n3292), .Z(n3342));
  OR2 U3252 ( .A(n3345), .B(n3346), .Z(n3335));
  IV2 U3253 ( .A(n3347), .Z(n3346));
  OR2 U3254 ( .A(n3348), .B(n3349), .Z(n3347));
  AN2 U3255 ( .A(n3349), .B(n3348), .Z(n3345));
  AN2 U3256 ( .A(n3350), .B(n3351), .Z(n3348));
  OR2 U3257 ( .A(n3352), .B(n3353), .Z(n3351));
  IV2 U3258 ( .A(n3354), .Z(n3353));
  OR2 U3259 ( .A(n3354), .B(n3355), .Z(n3350));
  OR2 U3260 ( .A(n3356), .B(n3357), .Z(n3354));
  OR2 U3261 ( .A(n3358), .B(n3359), .Z(n3357));
  AN2 U3262 ( .A(n3360), .B(n3361), .Z(n3359));
  AN2 U3263 ( .A(n3362), .B(n3363), .Z(n3360));
  OR2 U3264 ( .A(n3364), .B(n3365), .Z(n3362));
  OR2 U3265 ( .A(n3366), .B(n3367), .Z(n3365));
  AN2 U3266 ( .A(n3368), .B(n3369), .Z(n3367));
  AN2 U3267 ( .A(n3370), .B(n3371), .Z(n3368));
  AN2 U3268 ( .A(n3372), .B(n3373), .Z(n3366));
  AN2 U3269 ( .A(n3374), .B(n3375), .Z(n3372));
  OR2 U3270 ( .A(n3376), .B(n3377), .Z(n3374));
  OR2 U3271 ( .A(n3378), .B(n3379), .Z(n3377));
  AN2 U3272 ( .A(n2837), .B(n3380), .Z(n3379));
  AN2 U3273 ( .A(pi060), .B(n3381), .Z(n3378));
  AN2 U3274 ( .A(n3382), .B(n3369), .Z(n3364));
  AN2 U3275 ( .A(n3369), .B(n3383), .Z(n3358));
  OR2 U3276 ( .A(n3384), .B(n3385), .Z(n3383));
  OR2 U3277 ( .A(n3386), .B(n3387), .Z(n3385));
  AN2 U3278 ( .A(n3370), .B(n3388), .Z(n3387));
  OR2 U3279 ( .A(n3389), .B(n3390), .Z(n3388));
  AN2 U3280 ( .A(n3391), .B(n3392), .Z(n3390));
  AN2 U3281 ( .A(n3393), .B(n3394), .Z(n3386));
  OR2 U3282 ( .A(n3395), .B(n3396), .Z(n3394));
  OR2 U3283 ( .A(n3321), .B(n3397), .Z(n3396));
  AN2 U3284 ( .A(n3398), .B(n3399), .Z(n3397));
  AN2 U3285 ( .A(n3400), .B(n3401), .Z(n3395));
  OR2 U3286 ( .A(n3402), .B(n3371), .Z(n3400));
  AN2 U3287 ( .A(n3403), .B(n3404), .Z(n3402));
  AN2 U3288 ( .A(pi060), .B(po071), .Z(n3403));
  OR2 U3289 ( .A(n3405), .B(n3406), .Z(n3384));
  AN2 U3290 ( .A(n3407), .B(n3363), .Z(n3406));
  AN2 U3291 ( .A(n3408), .B(n3401), .Z(n3407));
  OR2 U3292 ( .A(n3409), .B(n3410), .Z(n3408));
  AN2 U3293 ( .A(n3411), .B(n3412), .Z(n3409));
  OR2 U3294 ( .A(n3413), .B(n3414), .Z(n3411));
  AN2 U3295 ( .A(n3415), .B(n3370), .Z(n3414));
  OR2 U3296 ( .A(n3416), .B(n3417), .Z(n3415));
  AN2 U3297 ( .A(n3418), .B(n3381), .Z(n3413));
  AN2 U3298 ( .A(n3393), .B(n3419), .Z(n3418));
  AN2 U3299 ( .A(n3420), .B(po027), .Z(n3405));
  OR2 U3300 ( .A(n3421), .B(n3422), .Z(n3420));
  OR2 U3301 ( .A(n3423), .B(n3424), .Z(n3422));
  AN2 U3302 ( .A(n3410), .B(n3361), .Z(n3424));
  IV2 U3303 ( .A(n3425), .Z(n3410));
  AN2 U3304 ( .A(n3426), .B(n3401), .Z(n3423));
  OR2 U3305 ( .A(n3427), .B(n3382), .Z(n3426));
  IV2 U3306 ( .A(n3428), .Z(n3382));
  OR2 U3307 ( .A(n3429), .B(n3430), .Z(n3421));
  AN2 U3308 ( .A(n3431), .B(n3370), .Z(n3430));
  AN2 U3309 ( .A(n3393), .B(n3432), .Z(n3429));
  OR2 U3310 ( .A(n3433), .B(n3434), .Z(n3432));
  AN2 U3311 ( .A(po071), .B(n3419), .Z(n3434));
  IV2 U3312 ( .A(n3435), .Z(n3369));
  OR2 U3313 ( .A(n3436), .B(n3375), .Z(n3435));
  AN2 U3314 ( .A(n3437), .B(n3438), .Z(n3436));
  AN2 U3315 ( .A(n3439), .B(n3440), .Z(n3438));
  OR2 U3316 ( .A(n3361), .B(n3441), .Z(n3440));
  AN2 U3317 ( .A(n3442), .B(n3443), .Z(n3441));
  OR2 U3318 ( .A(n3444), .B(n3445), .Z(n3443));
  OR2 U3319 ( .A(n3370), .B(n3446), .Z(n3445));
  OR2 U3320 ( .A(n3371), .B(n3380), .Z(n3444));
  AN2 U3321 ( .A(n3447), .B(n3448), .Z(n3442));
  OR2 U3322 ( .A(po027), .B(n3449), .Z(n3448));
  AN2 U3323 ( .A(n3450), .B(n3428), .Z(n3449));
  OR2 U3324 ( .A(n3371), .B(n3451), .Z(n3428));
  OR2 U3325 ( .A(n3370), .B(n3412), .Z(n3450));
  OR2 U3326 ( .A(n3363), .B(n3425), .Z(n3447));
  OR2 U3327 ( .A(n3427), .B(n3452), .Z(n3425));
  AN2 U3328 ( .A(n3453), .B(n3412), .Z(n3452));
  AN2 U3329 ( .A(n3371), .B(n3451), .Z(n3427));
  OR2 U3330 ( .A(n3401), .B(n3454), .Z(n3439));
  IV2 U3331 ( .A(n3455), .Z(n3454));
  AN2 U3332 ( .A(n3412), .B(n3456), .Z(n3455));
  OR2 U3333 ( .A(n3457), .B(n3458), .Z(n3456));
  AN2 U3334 ( .A(n3392), .B(n3393), .Z(n3458));
  AN2 U3335 ( .A(n3459), .B(n3460), .Z(n3437));
  OR2 U3336 ( .A(n3457), .B(n3461), .Z(n3460));
  AN2 U3337 ( .A(n3462), .B(n3463), .Z(n3459));
  OR2 U3338 ( .A(n3464), .B(n3370), .Z(n3463));
  IV2 U3339 ( .A(n3465), .Z(n3464));
  OR2 U3340 ( .A(n3389), .B(n3431), .Z(n3465));
  AN2 U3341 ( .A(n3466), .B(n3419), .Z(n3431));
  AN2 U3342 ( .A(n3467), .B(n3468), .Z(n3389));
  IV2 U3343 ( .A(n3469), .Z(n3468));
  OR2 U3344 ( .A(n3417), .B(n3470), .Z(n3469));
  AN2 U3345 ( .A(n3471), .B(n3399), .Z(n3470));
  OR2 U3346 ( .A(n3371), .B(n3446), .Z(n3471));
  OR2 U3347 ( .A(n3472), .B(n3393), .Z(n3462));
  AN2 U3348 ( .A(n3473), .B(n3474), .Z(n3472));
  AN2 U3349 ( .A(n3475), .B(n3476), .Z(n3474));
  OR2 U3350 ( .A(n3412), .B(n3477), .Z(n3476));
  AN2 U3351 ( .A(n3478), .B(n3261), .Z(n3475));
  IV2 U3352 ( .A(n3479), .Z(n3478));
  AN2 U3353 ( .A(n3361), .B(n3480), .Z(n3479));
  AN2 U3354 ( .A(n3481), .B(n3482), .Z(n3473));
  OR2 U3355 ( .A(n3483), .B(n3380), .Z(n3482));
  AN2 U3356 ( .A(n3484), .B(n3461), .Z(n3483));
  OR2 U3357 ( .A(n3371), .B(n3485), .Z(n3484));
  IV2 U3358 ( .A(n3433), .Z(n3481));
  OR2 U3359 ( .A(n3486), .B(n3417), .Z(n3433));
  AN2 U3360 ( .A(n3404), .B(n3381), .Z(n3417));
  AN2 U3361 ( .A(n3487), .B(n3380), .Z(n3486));
  AN2 U3362 ( .A(n3488), .B(n3375), .Z(n3356));
  OR2 U3363 ( .A(n3489), .B(n3490), .Z(n3375));
  AN2 U3364 ( .A(n3225), .B(n3491), .Z(n3489));
  OR2 U3365 ( .A(n3492), .B(n3493), .Z(n3491));
  AN2 U3366 ( .A(n3494), .B(n3495), .Z(n3492));
  OR2 U3367 ( .A(n3496), .B(n3497), .Z(n3488));
  OR2 U3368 ( .A(n3498), .B(n3499), .Z(n3497));
  AN2 U3369 ( .A(n3371), .B(n3500), .Z(n3499));
  OR2 U3370 ( .A(n3501), .B(n3502), .Z(n3500));
  OR2 U3371 ( .A(n3503), .B(n3504), .Z(n3502));
  AN2 U3372 ( .A(n3505), .B(n3401), .Z(n3504));
  OR2 U3373 ( .A(n3506), .B(n3507), .Z(n3505));
  AN2 U3374 ( .A(n3508), .B(n3509), .Z(n3507));
  OR2 U3375 ( .A(n3510), .B(n3511), .Z(n3509));
  OR2 U3376 ( .A(n3398), .B(n3487), .Z(n3511));
  AN2 U3377 ( .A(n3512), .B(n2837), .Z(n3487));
  AN2 U3378 ( .A(n3404), .B(pi060), .Z(n3510));
  AN2 U3379 ( .A(n3513), .B(po027), .Z(n3506));
  AN2 U3380 ( .A(n3514), .B(n3515), .Z(n3513));
  OR2 U3381 ( .A(n3516), .B(n3517), .Z(n3515));
  OR2 U3382 ( .A(n3321), .B(n3373), .Z(n3514));
  AN2 U3383 ( .A(n3518), .B(n3467), .Z(n3503));
  AN2 U3384 ( .A(n3404), .B(n3519), .Z(n3518));
  OR2 U3385 ( .A(n3520), .B(n3521), .Z(n3501));
  AN2 U3386 ( .A(n3522), .B(n3517), .Z(n3521));
  AN2 U3387 ( .A(n3516), .B(n3363), .Z(n3522));
  AN2 U3388 ( .A(n3373), .B(n3523), .Z(n3520));
  OR2 U3389 ( .A(n3524), .B(n3525), .Z(n3523));
  AN2 U3390 ( .A(n3361), .B(n3526), .Z(n3524));
  OR2 U3391 ( .A(n3527), .B(n3321), .Z(n3526));
  AN2 U3392 ( .A(n3519), .B(n3528), .Z(n3498));
  OR2 U3393 ( .A(n3529), .B(n3530), .Z(n3528));
  OR2 U3394 ( .A(n3392), .B(n3531), .Z(n3530));
  AN2 U3395 ( .A(n3376), .B(n3412), .Z(n3531));
  OR2 U3396 ( .A(n3532), .B(n3321), .Z(n3376));
  AN2 U3397 ( .A(n3533), .B(n3399), .Z(n3532));
  AN2 U3398 ( .A(n3534), .B(n3381), .Z(n3529));
  OR2 U3399 ( .A(n3535), .B(n3536), .Z(n3519));
  AN2 U3400 ( .A(n3537), .B(po027), .Z(n3536));
  AN2 U3401 ( .A(n3538), .B(n3363), .Z(n3535));
  AN2 U3402 ( .A(n3517), .B(n3401), .Z(n3538));
  OR2 U3403 ( .A(n3539), .B(n3540), .Z(n3496));
  AN2 U3404 ( .A(n3541), .B(n3542), .Z(n3540));
  OR2 U3405 ( .A(n3543), .B(n3544), .Z(n3542));
  AN2 U3406 ( .A(n3453), .B(po071), .Z(n3544));
  AN2 U3407 ( .A(n3480), .B(n3534), .Z(n3543));
  AN2 U3408 ( .A(n3545), .B(n3546), .Z(n3541));
  OR2 U3409 ( .A(n3361), .B(n3547), .Z(n3546));
  AN2 U3410 ( .A(n3508), .B(n3412), .Z(n3547));
  OR2 U3411 ( .A(n3401), .B(n3548), .Z(n3545));
  IV2 U3412 ( .A(n3508), .Z(n3548));
  OR2 U3413 ( .A(n3549), .B(n3550), .Z(n3508));
  AN2 U3414 ( .A(n3373), .B(n3363), .Z(n3550));
  AN2 U3415 ( .A(n3517), .B(po027), .Z(n3549));
  AN2 U3416 ( .A(n3551), .B(n3467), .Z(n3539));
  AN2 U3417 ( .A(n3552), .B(n3381), .Z(n3551));
  OR2 U3418 ( .A(n3553), .B(n3554), .Z(n3552));
  AN2 U3419 ( .A(n3537), .B(n3363), .Z(n3554));
  AN2 U3420 ( .A(n3555), .B(po027), .Z(n3553));
  IV2 U3421 ( .A(n3537), .Z(n3555));
  OR2 U3422 ( .A(n3556), .B(n3557), .Z(n3537));
  AN2 U3423 ( .A(n3373), .B(n3401), .Z(n3557));
  AN2 U3424 ( .A(n3517), .B(n3361), .Z(n3556));
  IV2 U3425 ( .A(n3373), .Z(n3517));
  OR2 U3426 ( .A(n3558), .B(n3559), .Z(n3373));
  AN2 U3427 ( .A(n3370), .B(n3560), .Z(n3559));
  OR2 U3428 ( .A(n3561), .B(n3562), .Z(n3560));
  OR2 U3429 ( .A(n3361), .B(n3563), .Z(n3562));
  AN2 U3430 ( .A(n3321), .B(po027), .Z(n3563));
  OR2 U3431 ( .A(n3564), .B(n3565), .Z(n3561));
  OR2 U3432 ( .A(n3527), .B(n3566), .Z(n3565));
  AN2 U3433 ( .A(po027), .B(n3398), .Z(n3527));
  AN2 U3434 ( .A(n3404), .B(n3567), .Z(n3564));
  AN2 U3435 ( .A(n3393), .B(n3568), .Z(n3558));
  OR2 U3436 ( .A(n3569), .B(n3570), .Z(n3568));
  AN2 U3437 ( .A(n3571), .B(n3401), .Z(n3570));
  OR2 U3438 ( .A(n3516), .B(n3572), .Z(n3571));
  AN2 U3439 ( .A(n3419), .B(n3363), .Z(n3572));
  AN2 U3440 ( .A(po104), .B(n3453), .Z(n3516));
  AN2 U3441 ( .A(n3573), .B(n3467), .Z(n3569));
  AN2 U3442 ( .A(n3261), .B(n3533), .Z(n3467));
  AN2 U3443 ( .A(n3404), .B(po027), .Z(n3573));
  OR2 U3444 ( .A(n3574), .B(n3575), .Z(n3349));
  AN2 U3445 ( .A(n3576), .B(n3247), .Z(n3575));
  IV2 U3446 ( .A(n3577), .Z(n3576));
  AN2 U3447 ( .A(n3225), .B(n3577), .Z(n3574));
  OR2 U3448 ( .A(n3578), .B(n3579), .Z(n3577));
  OR2 U3449 ( .A(n3580), .B(n3581), .Z(n3579));
  OR2 U3450 ( .A(n3582), .B(n3583), .Z(n3581));
  AN2 U3451 ( .A(n3584), .B(n2837), .Z(n3583));
  OR2 U3452 ( .A(n3585), .B(n3586), .Z(n3584));
  OR2 U3453 ( .A(n3587), .B(n3588), .Z(n3586));
  AN2 U3454 ( .A(n3589), .B(n3590), .Z(n3588));
  AN2 U3455 ( .A(n3591), .B(n3592), .Z(n3589));
  OR2 U3456 ( .A(n3593), .B(n3355), .Z(n3592));
  AN2 U3457 ( .A(n3594), .B(n3595), .Z(n3591));
  OR2 U3458 ( .A(n3596), .B(n3597), .Z(n3595));
  OR2 U3459 ( .A(pi003), .B(n3598), .Z(n3594));
  AN2 U3460 ( .A(n3599), .B(n3600), .Z(n3587));
  OR2 U3461 ( .A(n3601), .B(n3602), .Z(n3600));
  OR2 U3462 ( .A(n3603), .B(n3604), .Z(n3602));
  AN2 U3463 ( .A(n3605), .B(n3593), .Z(n3604));
  AN2 U3464 ( .A(n3606), .B(n3607), .Z(n3603));
  OR2 U3465 ( .A(n3608), .B(n3609), .Z(n3601));
  AN2 U3466 ( .A(n3610), .B(pi003), .Z(n3609));
  AN2 U3467 ( .A(n3611), .B(n3612), .Z(n3610));
  AN2 U3468 ( .A(n3613), .B(n3597), .Z(n3608));
  OR2 U3469 ( .A(n3614), .B(n3615), .Z(n3613));
  AN2 U3470 ( .A(n3598), .B(n3616), .Z(n3615));
  AN2 U3471 ( .A(n3617), .B(n3593), .Z(n3614));
  AN2 U3472 ( .A(n3618), .B(n3619), .Z(n3585));
  AN2 U3473 ( .A(n3620), .B(n3590), .Z(n3618));
  OR2 U3474 ( .A(n3621), .B(n3622), .Z(n3620));
  OR2 U3475 ( .A(n3494), .B(n3606), .Z(n3622));
  AN2 U3476 ( .A(pi003), .B(n3623), .Z(n3606));
  AN2 U3477 ( .A(n3616), .B(po011), .Z(n3623));
  AN2 U3478 ( .A(n3624), .B(n3625), .Z(n3621));
  AN2 U3479 ( .A(n3616), .B(n3597), .Z(n3624));
  AN2 U3480 ( .A(pi192), .B(n3626), .Z(n3582));
  OR2 U3481 ( .A(n3627), .B(n3628), .Z(n3626));
  OR2 U3482 ( .A(n3629), .B(n3630), .Z(n3628));
  AN2 U3483 ( .A(n3631), .B(n3632), .Z(n3630));
  AN2 U3484 ( .A(n3633), .B(n3634), .Z(n3631));
  OR2 U3485 ( .A(n3635), .B(n3355), .Z(n3634));
  AN2 U3486 ( .A(n3636), .B(n3637), .Z(n3633));
  OR2 U3487 ( .A(n3596), .B(n3638), .Z(n3637));
  AN2 U3488 ( .A(n3639), .B(n3339), .Z(n3596));
  OR2 U3489 ( .A(pi098), .B(n3598), .Z(n3636));
  AN2 U3490 ( .A(n3640), .B(n3641), .Z(n3629));
  OR2 U3491 ( .A(n3642), .B(n3643), .Z(n3641));
  OR2 U3492 ( .A(n3644), .B(n3645), .Z(n3643));
  AN2 U3493 ( .A(n3605), .B(n3635), .Z(n3645));
  OR2 U3494 ( .A(n3646), .B(n3647), .Z(n3605));
  AN2 U3495 ( .A(n3648), .B(n3493), .Z(n3647));
  AN2 U3496 ( .A(n3341), .B(n3639), .Z(n3646));
  AN2 U3497 ( .A(n3649), .B(n3607), .Z(n3644));
  OR2 U3498 ( .A(n3650), .B(n3651), .Z(n3642));
  AN2 U3499 ( .A(n3652), .B(pi098), .Z(n3651));
  AN2 U3500 ( .A(n3653), .B(n3612), .Z(n3652));
  AN2 U3501 ( .A(n3654), .B(n3638), .Z(n3650));
  OR2 U3502 ( .A(n3655), .B(n3656), .Z(n3654));
  AN2 U3503 ( .A(n3598), .B(n3657), .Z(n3656));
  OR2 U3504 ( .A(n3658), .B(n3659), .Z(n3598));
  AN2 U3505 ( .A(n3660), .B(n3493), .Z(n3659));
  AN2 U3506 ( .A(po011), .B(n3612), .Z(n3660));
  AN2 U3507 ( .A(n3625), .B(n3661), .Z(n3658));
  AN2 U3508 ( .A(n3617), .B(n3635), .Z(n3655));
  AN2 U3509 ( .A(n3625), .B(n3493), .Z(n3617));
  AN2 U3510 ( .A(n3662), .B(n3619), .Z(n3627));
  AN2 U3511 ( .A(n3663), .B(n3632), .Z(n3662));
  OR2 U3512 ( .A(n3664), .B(n3665), .Z(n3663));
  OR2 U3513 ( .A(n3494), .B(n3649), .Z(n3665));
  AN2 U3514 ( .A(pi098), .B(n3666), .Z(n3649));
  AN2 U3515 ( .A(n3657), .B(po011), .Z(n3666));
  AN2 U3516 ( .A(n3612), .B(n3667), .Z(n3494));
  AN2 U3517 ( .A(n3668), .B(n3625), .Z(n3664));
  AN2 U3518 ( .A(n3657), .B(n3638), .Z(n3668));
  OR2 U3519 ( .A(n3669), .B(n3670), .Z(n3580));
  AN2 U3520 ( .A(n3671), .B(po011), .Z(n3670));
  AN2 U3521 ( .A(n3672), .B(n3612), .Z(n3671));
  AN2 U3522 ( .A(n3673), .B(n3674), .Z(n3672));
  OR2 U3523 ( .A(pi192), .B(n3675), .Z(n3674));
  AN2 U3524 ( .A(n3676), .B(n3597), .Z(n3675));
  OR2 U3525 ( .A(n3677), .B(n3678), .Z(n3676));
  AN2 U3526 ( .A(n3679), .B(n3680), .Z(n3677));
  AN2 U3527 ( .A(n3599), .B(n3661), .Z(n3679));
  OR2 U3528 ( .A(n2837), .B(n3681), .Z(n3673));
  AN2 U3529 ( .A(n3682), .B(n3638), .Z(n3681));
  OR2 U3530 ( .A(n3683), .B(n3684), .Z(n3682));
  AN2 U3531 ( .A(n3685), .B(n3686), .Z(n3683));
  AN2 U3532 ( .A(n3640), .B(n3661), .Z(n3685));
  AN2 U3533 ( .A(n3687), .B(n3688), .Z(n3669));
  OR2 U3534 ( .A(n3689), .B(n3690), .Z(n3687));
  OR2 U3535 ( .A(n3691), .B(n3692), .Z(n3690));
  AN2 U3536 ( .A(n3693), .B(n3612), .Z(n3692));
  AN2 U3537 ( .A(n3619), .B(n3694), .Z(n3693));
  OR2 U3538 ( .A(n3695), .B(n3696), .Z(n3694));
  OR2 U3539 ( .A(n3697), .B(n3698), .Z(n3696));
  AN2 U3540 ( .A(n3699), .B(n3616), .Z(n3698));
  AN2 U3541 ( .A(n3700), .B(n3657), .Z(n3697));
  AN2 U3542 ( .A(n3341), .B(n3701), .Z(n3695));
  AN2 U3543 ( .A(n3493), .B(n3352), .Z(n3619));
  AN2 U3544 ( .A(n3625), .B(n3702), .Z(n3691));
  OR2 U3545 ( .A(n3703), .B(n3704), .Z(n3702));
  AN2 U3546 ( .A(n3705), .B(n3706), .Z(n3704));
  OR2 U3547 ( .A(n3684), .B(n3707), .Z(n3706));
  OR2 U3548 ( .A(n3708), .B(n3709), .Z(n3707));
  AN2 U3549 ( .A(n3710), .B(n3640), .Z(n3709));
  OR2 U3550 ( .A(n3711), .B(n3712), .Z(n3710));
  AN2 U3551 ( .A(n3607), .B(n3686), .Z(n3712));
  AN2 U3552 ( .A(n3493), .B(n3713), .Z(n3711));
  IV2 U3553 ( .A(n3686), .Z(n3713));
  AN2 U3554 ( .A(n3653), .B(n3632), .Z(n3708));
  OR2 U3555 ( .A(n3714), .B(n3715), .Z(n3653));
  AN2 U3556 ( .A(n3686), .B(n3493), .Z(n3714));
  AN2 U3557 ( .A(n3635), .B(n3339), .Z(n3686));
  AN2 U3558 ( .A(n3607), .B(n3716), .Z(n3684));
  AN2 U3559 ( .A(n3632), .B(n3657), .Z(n3716));
  AN2 U3560 ( .A(n3717), .B(n3718), .Z(n3703));
  OR2 U3561 ( .A(n3678), .B(n3719), .Z(n3718));
  OR2 U3562 ( .A(n3720), .B(n3721), .Z(n3719));
  AN2 U3563 ( .A(n3722), .B(n3599), .Z(n3721));
  OR2 U3564 ( .A(n3723), .B(n3724), .Z(n3722));
  AN2 U3565 ( .A(n3680), .B(n3607), .Z(n3724));
  AN2 U3566 ( .A(n3493), .B(n3725), .Z(n3723));
  IV2 U3567 ( .A(n3680), .Z(n3725));
  AN2 U3568 ( .A(n3611), .B(n3590), .Z(n3720));
  OR2 U3569 ( .A(n3726), .B(n3715), .Z(n3611));
  AN2 U3570 ( .A(n3341), .B(n3607), .Z(n3715));
  AN2 U3571 ( .A(n3680), .B(n3493), .Z(n3726));
  AN2 U3572 ( .A(n3593), .B(n3339), .Z(n3680));
  AN2 U3573 ( .A(n3607), .B(n3727), .Z(n3678));
  AN2 U3574 ( .A(n3590), .B(n3616), .Z(n3727));
  AN2 U3575 ( .A(n3661), .B(n3352), .Z(n3607));
  AN2 U3576 ( .A(n3639), .B(n3728), .Z(n3689));
  OR2 U3577 ( .A(n3729), .B(n3730), .Z(n3728));
  OR2 U3578 ( .A(n3731), .B(n3732), .Z(n3730));
  AN2 U3579 ( .A(n3733), .B(pi192), .Z(n3732));
  AN2 U3580 ( .A(n3640), .B(n3657), .Z(n3733));
  AN2 U3581 ( .A(n3734), .B(n2837), .Z(n3731));
  AN2 U3582 ( .A(n3599), .B(n3616), .Z(n3734));
  IV2 U3583 ( .A(n3590), .Z(n3599));
  AN2 U3584 ( .A(n3735), .B(n3355), .Z(n3729));
  OR2 U3585 ( .A(n3339), .B(n3736), .Z(n3735));
  OR2 U3586 ( .A(n3737), .B(n3738), .Z(n3578));
  AN2 U3587 ( .A(n3355), .B(n3739), .Z(n3738));
  OR2 U3588 ( .A(n3740), .B(n3741), .Z(n3739));
  AN2 U3589 ( .A(n3742), .B(n3625), .Z(n3741));
  AN2 U3590 ( .A(n3743), .B(n3744), .Z(n3742));
  OR2 U3591 ( .A(n3661), .B(n3688), .Z(n3744));
  OR2 U3592 ( .A(po011), .B(n3745), .Z(n3743));
  AN2 U3593 ( .A(n3493), .B(n3746), .Z(n3745));
  AN2 U3594 ( .A(n3747), .B(n3639), .Z(n3740));
  AN2 U3595 ( .A(n3661), .B(n3612), .Z(n3639));
  AN2 U3596 ( .A(n3736), .B(n3746), .Z(n3747));
  OR2 U3597 ( .A(n3292), .B(n3344), .Z(n3736));
  IV2 U3598 ( .A(n3291), .Z(n3292));
  AN2 U3599 ( .A(n3748), .B(n3648), .Z(n3737));
  OR2 U3600 ( .A(n3749), .B(n3750), .Z(n3648));
  AN2 U3601 ( .A(n3625), .B(po011), .Z(n3750));
  IV2 U3602 ( .A(n3612), .Z(n3625));
  AN2 U3603 ( .A(n3751), .B(n3688), .Z(n3749));
  AN2 U3604 ( .A(n3339), .B(n3612), .Z(n3751));
  OR2 U3605 ( .A(n3752), .B(n3753), .Z(n3612));
  OR2 U3606 ( .A(n3754), .B(n3755), .Z(n3753));
  AN2 U3607 ( .A(n3756), .B(n3757), .Z(n3755));
  OR2 U3608 ( .A(n3758), .B(n3759), .Z(n3752));
  AN2 U3609 ( .A(n3760), .B(n3761), .Z(n3759));
  AN2 U3610 ( .A(n3661), .B(n3762), .Z(n3748));
  OR2 U3611 ( .A(n3763), .B(n3764), .Z(po087));
  OR2 U3612 ( .A(po042), .B(n3765), .Z(n3764));
  OR2 U3613 ( .A(po029), .B(po022), .Z(n3765));
  OR2 U3614 ( .A(n3766), .B(n3767), .Z(n3763));
  OR2 U3615 ( .A(po080), .B(po056), .Z(n3767));
  OR2 U3616 ( .A(po105), .B(po083), .Z(n3766));
  IV2 U3617 ( .A(n3768), .Z(po105));
  AN2 U3618 ( .A(n3769), .B(n3770), .Z(n3768));
  AN2 U3619 ( .A(pi034), .B(pi007), .Z(n3770));
  AN2 U3620 ( .A(pi139), .B(pi120), .Z(n3769));
  OR2 U3621 ( .A(n3771), .B(n3772), .Z(po086));
  AN2 U3622 ( .A(n3773), .B(n3774), .Z(n3772));
  OR2 U3623 ( .A(n3775), .B(n3776), .Z(n3774));
  AN2 U3624 ( .A(n3777), .B(n3778), .Z(n3771));
  AN2 U3625 ( .A(n3779), .B(n3780), .Z(n3777));
  OR2 U3626 ( .A(po025), .B(n3781), .Z(n3779));
  IV2 U3627 ( .A(n3782), .Z(po083));
  AN2 U3628 ( .A(n3783), .B(n3784), .Z(n3782));
  AN2 U3629 ( .A(pi067), .B(pi041), .Z(n3784));
  AN2 U3630 ( .A(pi104), .B(pi070), .Z(n3783));
  OR2 U3631 ( .A(n3785), .B(n3786), .Z(po081));
  AN2 U3632 ( .A(n2862), .B(n3787), .Z(n3786));
  AN2 U3633 ( .A(n2930), .B(n3788), .Z(n3785));
  OR2 U3634 ( .A(n3146), .B(n3789), .Z(n3788));
  OR2 U3635 ( .A(n3790), .B(n3791), .Z(n3789));
  AN2 U3636 ( .A(n3792), .B(n2901), .Z(n3791));
  OR2 U3637 ( .A(n3793), .B(n3794), .Z(n3792));
  AN2 U3638 ( .A(pi192), .B(n2887), .Z(n3794));
  AN2 U3639 ( .A(n3795), .B(n2974), .Z(n3793));
  OR2 U3640 ( .A(n3796), .B(po031), .Z(n3795));
  AN2 U3641 ( .A(n2957), .B(n2837), .Z(n3796));
  AN2 U3642 ( .A(n3797), .B(n2935), .Z(n3790));
  AN2 U3643 ( .A(n2946), .B(n2837), .Z(n3797));
  OR2 U3644 ( .A(n3798), .B(n3799), .Z(po080));
  OR2 U3645 ( .A(n3800), .B(n3801), .Z(n3799));
  OR2 U3646 ( .A(n3802), .B(n3803), .Z(n3801));
  AN2 U3647 ( .A(n3804), .B(n2837), .Z(n3803));
  OR2 U3648 ( .A(n3805), .B(n3806), .Z(n3804));
  OR2 U3649 ( .A(n3807), .B(n3808), .Z(n3806));
  AN2 U3650 ( .A(n3809), .B(n3810), .Z(n3808));
  AN2 U3651 ( .A(n3811), .B(n3812), .Z(n3807));
  AN2 U3652 ( .A(n3813), .B(n3814), .Z(n3805));
  OR2 U3653 ( .A(n3815), .B(n3816), .Z(n3814));
  OR2 U3654 ( .A(n3817), .B(n3818), .Z(n3813));
  AN2 U3655 ( .A(pi192), .B(n3819), .Z(n3802));
  OR2 U3656 ( .A(n3820), .B(n3821), .Z(n3819));
  OR2 U3657 ( .A(n3822), .B(n3823), .Z(n3821));
  AN2 U3658 ( .A(n3824), .B(n3825), .Z(n3823));
  OR2 U3659 ( .A(n3826), .B(n3827), .Z(n3825));
  IV2 U3660 ( .A(n3828), .Z(n3824));
  AN2 U3661 ( .A(n3827), .B(n3826), .Z(n3828));
  OR2 U3662 ( .A(n3829), .B(n3830), .Z(n3826));
  AN2 U3663 ( .A(n3817), .B(n3171), .Z(n3830));
  AN2 U3664 ( .A(n3816), .B(pi033), .Z(n3829));
  IV2 U3665 ( .A(n3817), .Z(n3816));
  OR2 U3666 ( .A(n3831), .B(n3832), .Z(n3817));
  AN2 U3667 ( .A(n3833), .B(pi192), .Z(n3832));
  OR2 U3668 ( .A(n3834), .B(n3835), .Z(n3833));
  IV2 U3669 ( .A(n3836), .Z(n3835));
  OR2 U3670 ( .A(n3837), .B(n3838), .Z(n3836));
  AN2 U3671 ( .A(n3838), .B(n3837), .Z(n3834));
  AN2 U3672 ( .A(n3839), .B(n3840), .Z(n3837));
  OR2 U3673 ( .A(n3841), .B(pi013), .Z(n3840));
  IV2 U3674 ( .A(n3842), .Z(n3841));
  OR2 U3675 ( .A(n3843), .B(n3842), .Z(n3839));
  OR2 U3676 ( .A(n3844), .B(n3845), .Z(n3842));
  AN2 U3677 ( .A(pi026), .B(n3846), .Z(n3845));
  AN2 U3678 ( .A(pi077), .B(n3847), .Z(n3844));
  IV2 U3679 ( .A(pi013), .Z(n3843));
  OR2 U3680 ( .A(n3848), .B(n3849), .Z(n3838));
  AN2 U3681 ( .A(n3850), .B(n3136), .Z(n3849));
  AN2 U3682 ( .A(n3851), .B(pi088), .Z(n3848));
  IV2 U3683 ( .A(n3850), .Z(n3851));
  OR2 U3684 ( .A(n3852), .B(n3853), .Z(n3850));
  IV2 U3685 ( .A(n3854), .Z(n3853));
  OR2 U3686 ( .A(n3855), .B(pi157), .Z(n3854));
  AN2 U3687 ( .A(pi157), .B(n3855), .Z(n3852));
  IV2 U3688 ( .A(pi137), .Z(n3855));
  AN2 U3689 ( .A(n3856), .B(n3857), .Z(n3827));
  OR2 U3690 ( .A(n3858), .B(pi096), .Z(n3857));
  IV2 U3691 ( .A(n3859), .Z(n3858));
  OR2 U3692 ( .A(n3859), .B(n3199), .Z(n3856));
  OR2 U3693 ( .A(n3860), .B(n3861), .Z(n3859));
  AN2 U3694 ( .A(pi166), .B(n3862), .Z(n3861));
  IV2 U3695 ( .A(pi175), .Z(n3862));
  AN2 U3696 ( .A(pi175), .B(n3106), .Z(n3860));
  OR2 U3697 ( .A(n3863), .B(n3864), .Z(n3822));
  AN2 U3698 ( .A(n3865), .B(n3866), .Z(n3864));
  IV2 U3699 ( .A(n3867), .Z(n3863));
  OR2 U3700 ( .A(n3866), .B(n3865), .Z(n3867));
  OR2 U3701 ( .A(n3868), .B(n3869), .Z(n3865));
  AN2 U3702 ( .A(n3811), .B(n3870), .Z(n3869));
  IV2 U3703 ( .A(n3810), .Z(n3811));
  AN2 U3704 ( .A(pi016), .B(n3810), .Z(n3868));
  OR2 U3705 ( .A(n3871), .B(n3872), .Z(n3810));
  OR2 U3706 ( .A(n3873), .B(n3874), .Z(n3872));
  AN2 U3707 ( .A(n3875), .B(pi148), .Z(n3874));
  OR2 U3708 ( .A(n3876), .B(n3877), .Z(n3875));
  AN2 U3709 ( .A(n3878), .B(pi135), .Z(n3877));
  AN2 U3710 ( .A(n3879), .B(n3880), .Z(n3876));
  AN2 U3711 ( .A(n3881), .B(n3882), .Z(n3873));
  IV2 U3712 ( .A(pi148), .Z(n3882));
  OR2 U3713 ( .A(n3883), .B(n3884), .Z(n3881));
  AN2 U3714 ( .A(n3879), .B(pi135), .Z(n3884));
  OR2 U3715 ( .A(n3885), .B(n3886), .Z(n3879));
  AN2 U3716 ( .A(n3887), .B(n3888), .Z(n3886));
  AN2 U3717 ( .A(n3889), .B(n3890), .Z(n3885));
  AN2 U3718 ( .A(n3878), .B(n3880), .Z(n3883));
  OR2 U3719 ( .A(n3891), .B(n3892), .Z(n3878));
  AN2 U3720 ( .A(n3887), .B(n3890), .Z(n3892));
  AN2 U3721 ( .A(n3889), .B(n3888), .Z(n3891));
  IV2 U3722 ( .A(n3887), .Z(n3889));
  OR2 U3723 ( .A(n3893), .B(n3894), .Z(n3887));
  AN2 U3724 ( .A(n3895), .B(n3896), .Z(n3894));
  AN2 U3725 ( .A(n3897), .B(pi005), .Z(n3893));
  IV2 U3726 ( .A(n3895), .Z(n3897));
  OR2 U3727 ( .A(n3898), .B(n3899), .Z(n3895));
  AN2 U3728 ( .A(pi069), .B(n3900), .Z(n3899));
  IV2 U3729 ( .A(pi072), .Z(n3900));
  AN2 U3730 ( .A(pi072), .B(n3901), .Z(n3898));
  AN2 U3731 ( .A(n3902), .B(n3903), .Z(n3866));
  OR2 U3732 ( .A(n3904), .B(pi045), .Z(n3903));
  IV2 U3733 ( .A(n3905), .Z(n3902));
  AN2 U3734 ( .A(n3904), .B(pi045), .Z(n3905));
  AN2 U3735 ( .A(n3906), .B(n3907), .Z(n3904));
  OR2 U3736 ( .A(n3908), .B(pi158), .Z(n3907));
  OR2 U3737 ( .A(n3909), .B(pi079), .Z(n3906));
  OR2 U3738 ( .A(n3910), .B(n3911), .Z(n3820));
  AN2 U3739 ( .A(n3912), .B(n3913), .Z(n3911));
  AN2 U3740 ( .A(n3534), .B(n3914), .Z(n3912));
  AN2 U3741 ( .A(pi118), .B(n3915), .Z(n3910));
  OR2 U3742 ( .A(n3916), .B(n3917), .Z(n3915));
  AN2 U3743 ( .A(n3918), .B(pi060), .Z(n3917));
  AN2 U3744 ( .A(n3919), .B(n3534), .Z(n3916));
  AN2 U3745 ( .A(n3920), .B(n3921), .Z(n3919));
  AN2 U3746 ( .A(n3922), .B(n3923), .Z(n3800));
  OR2 U3747 ( .A(n3924), .B(n3925), .Z(n3923));
  OR2 U3748 ( .A(n3321), .B(n3926), .Z(n3925));
  AN2 U3749 ( .A(n3927), .B(n3928), .Z(n3924));
  AN2 U3750 ( .A(pi050), .B(pi118), .Z(n3928));
  AN2 U3751 ( .A(pi196), .B(n3534), .Z(n3927));
  OR2 U3752 ( .A(n3929), .B(n3930), .Z(n3798));
  OR2 U3753 ( .A(n3931), .B(n3932), .Z(n3930));
  AN2 U3754 ( .A(n3933), .B(n3533), .Z(n3932));
  AN2 U3755 ( .A(n3934), .B(n3913), .Z(n3933));
  OR2 U3756 ( .A(n3918), .B(n3935), .Z(n3934));
  OR2 U3757 ( .A(n3936), .B(n3937), .Z(n3935));
  AN2 U3758 ( .A(n3938), .B(n3921), .Z(n3937));
  AN2 U3759 ( .A(n3920), .B(n3261), .Z(n3938));
  AN2 U3760 ( .A(n3939), .B(n3922), .Z(n3936));
  AN2 U3761 ( .A(pi196), .B(n3940), .Z(n3939));
  AN2 U3762 ( .A(n3922), .B(n3941), .Z(n3918));
  AN2 U3763 ( .A(n3942), .B(n3943), .Z(n3941));
  AN2 U3764 ( .A(n3944), .B(n3945), .Z(n3931));
  AN2 U3765 ( .A(pi204), .B(n3946), .Z(n3944));
  IV2 U3766 ( .A(n3947), .Z(n3946));
  AN2 U3767 ( .A(n3948), .B(n3261), .Z(n3929));
  OR2 U3768 ( .A(n3949), .B(n3950), .Z(n3948));
  AN2 U3769 ( .A(n3947), .B(n3951), .Z(n3950));
  AN2 U3770 ( .A(n3952), .B(n3953), .Z(n3947));
  IV2 U3771 ( .A(n3954), .Z(n3953));
  AN2 U3772 ( .A(n3955), .B(n3956), .Z(n3954));
  OR2 U3773 ( .A(n3956), .B(n3955), .Z(n3952));
  OR2 U3774 ( .A(n3957), .B(n3958), .Z(n3955));
  AN2 U3775 ( .A(n3959), .B(n3960), .Z(n3958));
  IV2 U3776 ( .A(pi009), .Z(n3960));
  AN2 U3777 ( .A(pi009), .B(n3961), .Z(n3957));
  AN2 U3778 ( .A(n3962), .B(n3963), .Z(n3956));
  OR2 U3779 ( .A(n3964), .B(pi129), .Z(n3963));
  IV2 U3780 ( .A(n3965), .Z(n3964));
  OR2 U3781 ( .A(n3965), .B(n3966), .Z(n3962));
  OR2 U3782 ( .A(n3967), .B(n3968), .Z(n3965));
  AN2 U3783 ( .A(pi138), .B(n3969), .Z(n3968));
  AN2 U3784 ( .A(pi169), .B(n3970), .Z(n3967));
  IV2 U3785 ( .A(pi138), .Z(n3970));
  AN2 U3786 ( .A(n3971), .B(n3533), .Z(n3949));
  AN2 U3787 ( .A(n3914), .B(pi118), .Z(n3971));
  OR2 U3788 ( .A(n3972), .B(n3973), .Z(n3914));
  AN2 U3789 ( .A(n3920), .B(n3922), .Z(n3973));
  IV2 U3790 ( .A(n3921), .Z(n3922));
  AN2 U3791 ( .A(n3921), .B(n3974), .Z(n3972));
  IV2 U3792 ( .A(n3920), .Z(n3974));
  OR2 U3793 ( .A(n3975), .B(n3976), .Z(n3920));
  AN2 U3794 ( .A(pi050), .B(n3942), .Z(n3976));
  AN2 U3795 ( .A(pi196), .B(n3943), .Z(n3975));
  OR2 U3796 ( .A(n3977), .B(n3978), .Z(n3921));
  AN2 U3797 ( .A(n3979), .B(pi192), .Z(n3978));
  OR2 U3798 ( .A(n3980), .B(n3981), .Z(n3979));
  AN2 U3799 ( .A(n3982), .B(n3983), .Z(n3981));
  IV2 U3800 ( .A(n3984), .Z(n3980));
  OR2 U3801 ( .A(n3983), .B(n3982), .Z(n3984));
  OR2 U3802 ( .A(n3985), .B(n3986), .Z(n3982));
  IV2 U3803 ( .A(n3987), .Z(n3986));
  OR2 U3804 ( .A(n3988), .B(n3989), .Z(n3987));
  AN2 U3805 ( .A(n3988), .B(n3989), .Z(n3985));
  AN2 U3806 ( .A(n3990), .B(n3991), .Z(n3988));
  OR2 U3807 ( .A(n3992), .B(pi039), .Z(n3991));
  OR2 U3808 ( .A(n3993), .B(pi004), .Z(n3990));
  IV2 U3809 ( .A(pi039), .Z(n3993));
  AN2 U3810 ( .A(n3994), .B(n3995), .Z(n3983));
  OR2 U3811 ( .A(n3996), .B(pi068), .Z(n3995));
  IV2 U3812 ( .A(n3997), .Z(n3996));
  OR2 U3813 ( .A(n3997), .B(n3998), .Z(n3994));
  OR2 U3814 ( .A(n3999), .B(n4000), .Z(n3997));
  AN2 U3815 ( .A(pi098), .B(n4001), .Z(n4000));
  AN2 U3816 ( .A(pi171), .B(n3638), .Z(n3999));
  OR2 U3817 ( .A(pi037), .B(pi043), .Z(po078));
  OR2 U3818 ( .A(n4002), .B(n4003), .Z(po077));
  AN2 U3819 ( .A(n4004), .B(n4005), .Z(n4003));
  AN2 U3820 ( .A(n4006), .B(n4007), .Z(n4002));
  OR2 U3821 ( .A(n4008), .B(n4009), .Z(n4007));
  IV2 U3822 ( .A(pi090), .Z(po076));
  OR2 U3823 ( .A(n4010), .B(n4011), .Z(po075));
  AN2 U3824 ( .A(n4012), .B(n4013), .Z(n4011));
  OR2 U3825 ( .A(n4014), .B(n4015), .Z(n4012));
  OR2 U3826 ( .A(n4016), .B(n4017), .Z(n4015));
  OR2 U3827 ( .A(n4018), .B(n4019), .Z(n4014));
  AN2 U3828 ( .A(n4020), .B(n3314), .Z(n4019));
  OR2 U3829 ( .A(n4021), .B(n4022), .Z(n4020));
  AN2 U3830 ( .A(n3926), .B(n3328), .Z(n4022));
  OR2 U3831 ( .A(n3265), .B(n3326), .Z(n3328));
  AN2 U3832 ( .A(n4023), .B(pi204), .Z(n4021));
  AN2 U3833 ( .A(n3312), .B(n3261), .Z(n4023));
  OR2 U3834 ( .A(n4024), .B(n4025), .Z(n3312));
  AN2 U3835 ( .A(n3326), .B(n4026), .Z(n4024));
  AN2 U3836 ( .A(n4027), .B(n3320), .Z(n4018));
  OR2 U3837 ( .A(n4028), .B(n3321), .Z(n4027));
  AN2 U3838 ( .A(po040), .B(n4029), .Z(n4010));
  OR2 U3839 ( .A(n4030), .B(n4031), .Z(n4029));
  OR2 U3840 ( .A(n4032), .B(n4033), .Z(n4031));
  AN2 U3841 ( .A(n4034), .B(n3261), .Z(n4032));
  OR2 U3842 ( .A(n4035), .B(n4036), .Z(n4034));
  OR2 U3843 ( .A(n4037), .B(n4038), .Z(n4036));
  AN2 U3844 ( .A(n4039), .B(n3951), .Z(n4038));
  AN2 U3845 ( .A(n4025), .B(n3314), .Z(n4039));
  AN2 U3846 ( .A(n4040), .B(n4041), .Z(n4037));
  AN2 U3847 ( .A(n4042), .B(n3320), .Z(n4035));
  OR2 U3848 ( .A(n4043), .B(n4044), .Z(n4042));
  AN2 U3849 ( .A(pi204), .B(n4045), .Z(n4044));
  AN2 U3850 ( .A(n4046), .B(n4041), .Z(n4043));
  OR2 U3851 ( .A(n4047), .B(n4048), .Z(n4030));
  AN2 U3852 ( .A(n4049), .B(n4050), .Z(n4048));
  OR2 U3853 ( .A(n4051), .B(n4052), .Z(n4050));
  AN2 U3854 ( .A(n3321), .B(n3265), .Z(n4052));
  AN2 U3855 ( .A(n3951), .B(n4053), .Z(n4051));
  AN2 U3856 ( .A(n3326), .B(n3314), .Z(n4049));
  AN2 U3857 ( .A(n4054), .B(n4055), .Z(n4047));
  AN2 U3858 ( .A(n4056), .B(n4057), .Z(n4055));
  AN2 U3859 ( .A(n3945), .B(pi204), .Z(n4054));
  OR2 U3860 ( .A(n4058), .B(n4059), .Z(po073));
  AN2 U3861 ( .A(n4060), .B(n4061), .Z(n4059));
  AN2 U3862 ( .A(n3457), .B(n4062), .Z(n4058));
  OR2 U3863 ( .A(n4063), .B(n4064), .Z(po068));
  AN2 U3864 ( .A(n4065), .B(n4066), .Z(n4064));
  OR2 U3865 ( .A(n4067), .B(n4068), .Z(n4065));
  OR2 U3866 ( .A(n4069), .B(n4070), .Z(n4068));
  AN2 U3867 ( .A(n4071), .B(n4072), .Z(n4070));
  OR2 U3868 ( .A(n4073), .B(po059), .Z(n4071));
  AN2 U3869 ( .A(n4074), .B(n2837), .Z(n4073));
  AN2 U3870 ( .A(n4075), .B(n4076), .Z(n4069));
  AN2 U3871 ( .A(n3780), .B(n4077), .Z(n4075));
  AN2 U3872 ( .A(n4078), .B(n4079), .Z(n4063));
  OR2 U3873 ( .A(n4080), .B(n4081), .Z(n4079));
  OR2 U3874 ( .A(n4082), .B(n4083), .Z(n4081));
  AN2 U3875 ( .A(n4084), .B(n2837), .Z(n4083));
  AN2 U3876 ( .A(n4085), .B(pi192), .Z(n4082));
  AN2 U3877 ( .A(n3778), .B(n3776), .Z(n4080));
  OR2 U3878 ( .A(n4086), .B(n4087), .Z(n3776));
  OR2 U3879 ( .A(n4088), .B(n4089), .Z(po061));
  AN2 U3880 ( .A(n2861), .B(n4090), .Z(n4089));
  OR2 U3881 ( .A(n4091), .B(n4092), .Z(n4090));
  OR2 U3882 ( .A(n4093), .B(n4094), .Z(n4092));
  AN2 U3883 ( .A(n4095), .B(n2901), .Z(n4094));
  AN2 U3884 ( .A(n2862), .B(n2990), .Z(n4093));
  OR2 U3885 ( .A(n4096), .B(n4097), .Z(n4091));
  AN2 U3886 ( .A(n2880), .B(n4098), .Z(n4097));
  AN2 U3887 ( .A(n4099), .B(n4100), .Z(n4096));
  OR2 U3888 ( .A(n4101), .B(n4102), .Z(n4100));
  OR2 U3889 ( .A(n2978), .B(n4103), .Z(n4102));
  AN2 U3890 ( .A(n3222), .B(n2957), .Z(n4103));
  AN2 U3891 ( .A(n2935), .B(po031), .Z(n4101));
  IV2 U3892 ( .A(n2938), .Z(n2935));
  AN2 U3893 ( .A(n4104), .B(n2998), .Z(n4088));
  OR2 U3894 ( .A(n4105), .B(n4106), .Z(n4104));
  OR2 U3895 ( .A(n4107), .B(n4108), .Z(n4106));
  AN2 U3896 ( .A(n2892), .B(pi192), .Z(n4108));
  AN2 U3897 ( .A(n2929), .B(n2837), .Z(n4107));
  AN2 U3898 ( .A(n2930), .B(n3787), .Z(n4105));
  OR2 U3899 ( .A(n4109), .B(n4110), .Z(n3787));
  OR2 U3900 ( .A(n4111), .B(n4112), .Z(n4110));
  AN2 U3901 ( .A(n4113), .B(n2837), .Z(n4112));
  AN2 U3902 ( .A(n2876), .B(pi192), .Z(n4111));
  AN2 U3903 ( .A(pi200), .B(n4114), .Z(n4109));
  OR2 U3904 ( .A(n4115), .B(n2999), .Z(n4114));
  OR2 U3905 ( .A(n4116), .B(n4117), .Z(n2999));
  AN2 U3906 ( .A(n2938), .B(n2962), .Z(n4117));
  AN2 U3907 ( .A(pi192), .B(n2878), .Z(n4116));
  AN2 U3908 ( .A(n2918), .B(n2837), .Z(n4115));
  AN2 U3909 ( .A(n2938), .B(pi082), .Z(n2918));
  OR2 U3910 ( .A(n4118), .B(n4119), .Z(po060));
  OR2 U3911 ( .A(n4120), .B(n4121), .Z(n4119));
  AN2 U3912 ( .A(n4122), .B(n4123), .Z(n4121));
  OR2 U3913 ( .A(n4124), .B(n4125), .Z(n4123));
  AN2 U3914 ( .A(n4126), .B(n4127), .Z(n4124));
  OR2 U3915 ( .A(n4128), .B(n4129), .Z(n4126));
  AN2 U3916 ( .A(n4130), .B(n4131), .Z(n4122));
  OR2 U3917 ( .A(n4132), .B(n4133), .Z(n4131));
  AN2 U3918 ( .A(pi052), .B(n4134), .Z(n4132));
  OR2 U3919 ( .A(po064), .B(n4135), .Z(n4130));
  AN2 U3920 ( .A(n4136), .B(n4137), .Z(n4120));
  OR2 U3921 ( .A(n4138), .B(n4139), .Z(n4137));
  AN2 U3922 ( .A(n4140), .B(n4141), .Z(n4139));
  OR2 U3923 ( .A(n4142), .B(n4143), .Z(n4140));
  OR2 U3924 ( .A(n4144), .B(n4145), .Z(n4143));
  AN2 U3925 ( .A(po040), .B(n3321), .Z(n4145));
  AN2 U3926 ( .A(po103), .B(n4146), .Z(n4144));
  OR2 U3927 ( .A(n4147), .B(n3321), .Z(n4146));
  AN2 U3928 ( .A(n4148), .B(n4149), .Z(n4147));
  OR2 U3929 ( .A(po004), .B(n4150), .Z(n4149));
  OR2 U3930 ( .A(n4151), .B(n4152), .Z(n4142));
  OR2 U3931 ( .A(n4153), .B(n4154), .Z(n4152));
  IV2 U3932 ( .A(n4155), .Z(n4154));
  OR2 U3933 ( .A(n4156), .B(n4157), .Z(n4155));
  AN2 U3934 ( .A(n4158), .B(n4159), .Z(n4153));
  AN2 U3935 ( .A(n4160), .B(po004), .Z(n4151));
  AN2 U3936 ( .A(n3951), .B(po040), .Z(n4160));
  AN2 U3937 ( .A(po004), .B(n4161), .Z(n4138));
  AN2 U3938 ( .A(n4162), .B(n4163), .Z(n4136));
  OR2 U3939 ( .A(n4164), .B(n4134), .Z(n4163));
  AN2 U3940 ( .A(n4165), .B(po064), .Z(n4164));
  IV2 U3941 ( .A(n4166), .Z(n4165));
  OR2 U3942 ( .A(n4167), .B(n4125), .Z(n4166));
  OR2 U3943 ( .A(n4135), .B(n4168), .Z(n4162));
  OR2 U3944 ( .A(n4169), .B(n4170), .Z(n4168));
  AN2 U3945 ( .A(pi054), .B(n4167), .Z(n4170));
  AN2 U3946 ( .A(n4171), .B(n4133), .Z(n4169));
  IV2 U3947 ( .A(n4172), .Z(n4171));
  OR2 U3948 ( .A(n4173), .B(n4174), .Z(n4118));
  AN2 U3949 ( .A(n4175), .B(pi054), .Z(n4174));
  AN2 U3950 ( .A(n4176), .B(n4177), .Z(n4175));
  OR2 U3951 ( .A(n4178), .B(n4179), .Z(n4176));
  AN2 U3952 ( .A(n4134), .B(n4133), .Z(n4179));
  AN2 U3953 ( .A(n4135), .B(po064), .Z(n4178));
  AN2 U3954 ( .A(n4180), .B(n4135), .Z(n4173));
  IV2 U3955 ( .A(n4134), .Z(n4135));
  OR2 U3956 ( .A(n4181), .B(n4182), .Z(n4134));
  AN2 U3957 ( .A(n4183), .B(n4184), .Z(n4182));
  OR2 U3958 ( .A(n4185), .B(n4186), .Z(n4183));
  AN2 U3959 ( .A(n4187), .B(n4188), .Z(n4186));
  IV2 U3960 ( .A(n4189), .Z(n4188));
  OR2 U3961 ( .A(n4190), .B(n4191), .Z(n4187));
  AN2 U3962 ( .A(n4192), .B(n4193), .Z(n4191));
  OR2 U3963 ( .A(n4194), .B(n4195), .Z(n4193));
  AN2 U3964 ( .A(n4196), .B(n3261), .Z(n4195));
  OR2 U3965 ( .A(n4197), .B(n4198), .Z(n4196));
  AN2 U3966 ( .A(n4199), .B(po103), .Z(n4198));
  AN2 U3967 ( .A(n4200), .B(n4201), .Z(n4199));
  AN2 U3968 ( .A(n4202), .B(n4025), .Z(n4197));
  AN2 U3969 ( .A(n4203), .B(po091), .Z(n4202));
  AN2 U3970 ( .A(n4204), .B(n4205), .Z(n4190));
  OR2 U3971 ( .A(n3317), .B(n4206), .Z(n4204));
  OR2 U3972 ( .A(n4207), .B(n4208), .Z(n4206));
  AN2 U3973 ( .A(n4209), .B(n3314), .Z(n4208));
  IV2 U3974 ( .A(n4210), .Z(n4209));
  AN2 U3975 ( .A(n4210), .B(n4057), .Z(n4207));
  AN2 U3976 ( .A(po103), .B(n4148), .Z(n4210));
  AN2 U3977 ( .A(n4189), .B(n4211), .Z(n4185));
  OR2 U3978 ( .A(n4212), .B(n4213), .Z(n4211));
  AN2 U3979 ( .A(n4214), .B(n4205), .Z(n4213));
  OR2 U3980 ( .A(n3325), .B(n4215), .Z(n4214));
  OR2 U3981 ( .A(n4216), .B(n3329), .Z(n4215));
  AN2 U3982 ( .A(n4040), .B(n4217), .Z(n3329));
  AN2 U3983 ( .A(n4192), .B(n4218), .Z(n4212));
  OR2 U3984 ( .A(n4219), .B(n4220), .Z(n4218));
  OR2 U3985 ( .A(n4221), .B(n4222), .Z(n4220));
  AN2 U3986 ( .A(n4025), .B(n4201), .Z(n4222));
  IV2 U3987 ( .A(n4223), .Z(n4025));
  AN2 U3988 ( .A(po091), .B(n4200), .Z(n4221));
  OR2 U3989 ( .A(n4224), .B(n4225), .Z(n4189));
  AN2 U3990 ( .A(n4226), .B(n4227), .Z(n4225));
  IV2 U3991 ( .A(n4228), .Z(n4224));
  OR2 U3992 ( .A(n4227), .B(n4226), .Z(n4228));
  AN2 U3993 ( .A(n4229), .B(n4230), .Z(n4181));
  OR2 U3994 ( .A(n4231), .B(n4232), .Z(n4230));
  OR2 U3995 ( .A(n4233), .B(n4234), .Z(n4232));
  AN2 U3996 ( .A(n4235), .B(n4236), .Z(n4234));
  OR2 U3997 ( .A(n4237), .B(n4238), .Z(n4235));
  AN2 U3998 ( .A(n4239), .B(n4240), .Z(n4238));
  OR2 U3999 ( .A(n3325), .B(n4216), .Z(n4240));
  AN2 U4000 ( .A(po103), .B(n4194), .Z(n4216));
  AN2 U4001 ( .A(n3265), .B(n4040), .Z(n3325));
  AN2 U4002 ( .A(n4241), .B(n4242), .Z(n4237));
  OR2 U4003 ( .A(n4243), .B(n4219), .Z(n4241));
  OR2 U4004 ( .A(n4244), .B(n3321), .Z(n4219));
  AN2 U4005 ( .A(n4203), .B(n4223), .Z(n4244));
  AN2 U4006 ( .A(n4245), .B(n3314), .Z(n4243));
  OR2 U4007 ( .A(n4246), .B(po091), .Z(n4245));
  AN2 U4008 ( .A(n4247), .B(n3265), .Z(n4246));
  AN2 U4009 ( .A(n4248), .B(n4249), .Z(n4233));
  OR2 U4010 ( .A(n4250), .B(n4251), .Z(n4249));
  OR2 U4011 ( .A(n4252), .B(n4253), .Z(n4251));
  AN2 U4012 ( .A(po103), .B(n4254), .Z(n4253));
  OR2 U4013 ( .A(n4255), .B(n3330), .Z(n4254));
  AN2 U4014 ( .A(n3311), .B(n4242), .Z(n4255));
  AN2 U4015 ( .A(n4194), .B(n3265), .Z(n4252));
  AN2 U4016 ( .A(n4148), .B(n3311), .Z(n4194));
  AN2 U4017 ( .A(n4239), .B(n4256), .Z(n4250));
  OR2 U4018 ( .A(n4257), .B(n4258), .Z(n4256));
  OR2 U4019 ( .A(n3926), .B(n4259), .Z(n4258));
  AN2 U4020 ( .A(n4260), .B(n3314), .Z(n4259));
  OR2 U4021 ( .A(n4261), .B(n4262), .Z(n4257));
  AN2 U4022 ( .A(pi058), .B(pi129), .Z(n4262));
  AN2 U4023 ( .A(n4056), .B(n3966), .Z(n4261));
  AN2 U4024 ( .A(n4263), .B(n4264), .Z(n4231));
  AN2 U4025 ( .A(n4265), .B(n4266), .Z(n4264));
  OR2 U4026 ( .A(n4267), .B(n4236), .Z(n4266));
  AN2 U4027 ( .A(n4268), .B(pi058), .Z(n4267));
  AN2 U4028 ( .A(n4242), .B(n3265), .Z(n4268));
  OR2 U4029 ( .A(n4269), .B(n4248), .Z(n4265));
  IV2 U4030 ( .A(n4236), .Z(n4248));
  AN2 U4031 ( .A(n4270), .B(n4271), .Z(n4236));
  IV2 U4032 ( .A(n4272), .Z(n4271));
  AN2 U4033 ( .A(n4226), .B(n4141), .Z(n4272));
  OR2 U4034 ( .A(n4226), .B(n4141), .Z(n4270));
  OR2 U4035 ( .A(n4273), .B(n4274), .Z(n4226));
  IV2 U4036 ( .A(n4275), .Z(n4274));
  OR2 U4037 ( .A(n4276), .B(n4277), .Z(n4275));
  AN2 U4038 ( .A(n4277), .B(n4276), .Z(n4273));
  AN2 U4039 ( .A(n4278), .B(n4279), .Z(n4276));
  OR2 U4040 ( .A(n4280), .B(n4281), .Z(n4279));
  IV2 U4041 ( .A(n4282), .Z(n4280));
  OR2 U4042 ( .A(n4283), .B(n4282), .Z(n4278));
  OR2 U4043 ( .A(n4284), .B(n4285), .Z(n4282));
  AN2 U4044 ( .A(po040), .B(n4286), .Z(n4285));
  OR2 U4045 ( .A(n4017), .B(n4287), .Z(n4286));
  OR2 U4046 ( .A(n4288), .B(n4289), .Z(n4287));
  AN2 U4047 ( .A(n4290), .B(n3314), .Z(n4289));
  OR2 U4048 ( .A(n4291), .B(n3321), .Z(n4290));
  IV2 U4049 ( .A(n4292), .Z(n4288));
  OR2 U4050 ( .A(n4293), .B(n3314), .Z(n4292));
  OR2 U4051 ( .A(n4294), .B(n3330), .Z(n4017));
  AN2 U4052 ( .A(n4201), .B(n3926), .Z(n3330));
  AN2 U4053 ( .A(n3311), .B(pi204), .Z(n4294));
  AN2 U4054 ( .A(n4295), .B(n4013), .Z(n4284));
  OR2 U4055 ( .A(n4033), .B(n4296), .Z(n4295));
  OR2 U4056 ( .A(n4297), .B(n4298), .Z(n4296));
  AN2 U4057 ( .A(n4299), .B(n3314), .Z(n4298));
  AN2 U4058 ( .A(n4300), .B(n3261), .Z(n4299));
  OR2 U4059 ( .A(n4301), .B(n4302), .Z(n4300));
  AN2 U4060 ( .A(pi204), .B(n4203), .Z(n4302));
  AN2 U4061 ( .A(po091), .B(n4041), .Z(n4301));
  AN2 U4062 ( .A(n4040), .B(n4293), .Z(n4297));
  AN2 U4063 ( .A(n3311), .B(n3951), .Z(n4033));
  IV2 U4064 ( .A(n4260), .Z(n3311));
  OR2 U4065 ( .A(n3321), .B(n4057), .Z(n4260));
  IV2 U4066 ( .A(n4281), .Z(n4283));
  OR2 U4067 ( .A(n4303), .B(n4304), .Z(n4281));
  AN2 U4068 ( .A(n4305), .B(n4306), .Z(n4304));
  AN2 U4069 ( .A(n4307), .B(n3261), .Z(n4305));
  OR2 U4070 ( .A(n4308), .B(n4309), .Z(n4307));
  AN2 U4071 ( .A(pi065), .B(n4148), .Z(n4309));
  AN2 U4072 ( .A(n4310), .B(pi058), .Z(n4308));
  AN2 U4073 ( .A(n4311), .B(n4312), .Z(n4303));
  OR2 U4074 ( .A(n3961), .B(n4313), .Z(n4311));
  IV2 U4075 ( .A(n3959), .Z(n3961));
  OR2 U4076 ( .A(n4314), .B(n4315), .Z(n3959));
  AN2 U4077 ( .A(pi058), .B(n4150), .Z(n4315));
  AN2 U4078 ( .A(pi065), .B(n4316), .Z(n4314));
  OR2 U4079 ( .A(n4317), .B(n4318), .Z(n4277));
  AN2 U4080 ( .A(po004), .B(n3265), .Z(n4318));
  AN2 U4081 ( .A(po103), .B(n4319), .Z(n4317));
  AN2 U4082 ( .A(n4239), .B(pi058), .Z(n4269));
  AN2 U4083 ( .A(n4040), .B(n3261), .Z(n4263));
  AN2 U4084 ( .A(n4320), .B(n4167), .Z(n4180));
  OR2 U4085 ( .A(n4129), .B(n4127), .Z(n4320));
  AN2 U4086 ( .A(po023), .B(pi183), .Z(po058));
  IV2 U4087 ( .A(n4321), .Z(po056));
  AN2 U4088 ( .A(n4322), .B(n4323), .Z(n4321));
  AN2 U4089 ( .A(pi063), .B(pi010), .Z(n4323));
  AN2 U4090 ( .A(pi203), .B(pi073), .Z(n4322));
  OR2 U4091 ( .A(n4324), .B(n4325), .Z(po055));
  AN2 U4092 ( .A(n3015), .B(n4326), .Z(n4325));
  AN2 U4093 ( .A(n3018), .B(n4327), .Z(n4324));
  AN2 U4094 ( .A(n4328), .B(n4329), .Z(po053));
  OR2 U4095 ( .A(n4306), .B(n4330), .Z(n4329));
  IV2 U4096 ( .A(n4312), .Z(n4306));
  OR2 U4097 ( .A(n4331), .B(n4312), .Z(n4328));
  AN2 U4098 ( .A(n4332), .B(n3780), .Z(po051));
  OR2 U4099 ( .A(n4333), .B(n4334), .Z(n4332));
  OR2 U4100 ( .A(n4335), .B(n4336), .Z(po050));
  AN2 U4101 ( .A(n4337), .B(n4338), .Z(n4336));
  OR2 U4102 ( .A(n4339), .B(n4340), .Z(n4338));
  AN2 U4103 ( .A(n4087), .B(n4341), .Z(n4339));
  AN2 U4104 ( .A(n4342), .B(n4343), .Z(n4335));
  OR2 U4105 ( .A(n4344), .B(n4345), .Z(n4343));
  OR2 U4106 ( .A(n4346), .B(n4347), .Z(n4345));
  AN2 U4107 ( .A(n4067), .B(n4348), .Z(n4346));
  OR2 U4108 ( .A(n4349), .B(n4350), .Z(n4067));
  AN2 U4109 ( .A(n4351), .B(pi192), .Z(n4350));
  AN2 U4110 ( .A(n4072), .B(n3880), .Z(n4351));
  AN2 U4111 ( .A(n4352), .B(n3890), .Z(n4349));
  AN2 U4112 ( .A(n4353), .B(n3780), .Z(n4352));
  OR2 U4113 ( .A(n4354), .B(n4355), .Z(n4344));
  AN2 U4114 ( .A(n4356), .B(n3780), .Z(n4355));
  AN2 U4115 ( .A(n4357), .B(n4076), .Z(n4354));
  AN2 U4116 ( .A(n4072), .B(n4358), .Z(n4357));
  OR2 U4117 ( .A(n4359), .B(n4360), .Z(po049));
  AN2 U4118 ( .A(n3361), .B(n4361), .Z(n4360));
  OR2 U4119 ( .A(n4362), .B(n4363), .Z(n4361));
  AN2 U4120 ( .A(n4364), .B(n3451), .Z(n4362));
  IV2 U4121 ( .A(n3401), .Z(n3361));
  AN2 U4122 ( .A(n4365), .B(n3401), .Z(n4359));
  OR2 U4123 ( .A(n4366), .B(n4367), .Z(n4365));
  AN2 U4124 ( .A(n3453), .B(n4368), .Z(n4366));
  OR2 U4125 ( .A(n4369), .B(n3253), .Z(po048));
  AN2 U4126 ( .A(n4370), .B(n3255), .Z(n4369));
  OR2 U4127 ( .A(n4371), .B(n4372), .Z(n4370));
  AN2 U4128 ( .A(n4373), .B(n3259), .Z(n4371));
  AN2 U4129 ( .A(n4374), .B(n4242), .Z(n4373));
  OR2 U4130 ( .A(n4375), .B(n4376), .Z(po047));
  OR2 U4131 ( .A(n4377), .B(n4378), .Z(n4376));
  AN2 U4132 ( .A(n4379), .B(n4380), .Z(n4378));
  AN2 U4133 ( .A(n4381), .B(n3259), .Z(n4377));
  AN2 U4134 ( .A(n4382), .B(n4383), .Z(n4381));
  OR2 U4135 ( .A(po004), .B(n4384), .Z(n4383));
  OR2 U4136 ( .A(n3926), .B(n4385), .Z(n4384));
  AN2 U4137 ( .A(n4386), .B(pi065), .Z(n4385));
  AN2 U4138 ( .A(n4387), .B(n4157), .Z(n4386));
  OR2 U4139 ( .A(n4319), .B(n4388), .Z(n4382));
  OR2 U4140 ( .A(n4389), .B(n4390), .Z(n4388));
  AN2 U4141 ( .A(n4391), .B(n3321), .Z(n4390));
  AN2 U4142 ( .A(n4392), .B(n4310), .Z(n4389));
  AN2 U4143 ( .A(pi204), .B(n4387), .Z(n4392));
  OR2 U4144 ( .A(n4393), .B(n4394), .Z(n4375));
  AN2 U4145 ( .A(n4395), .B(n4319), .Z(n4394));
  OR2 U4146 ( .A(n4396), .B(n4397), .Z(n4395));
  AN2 U4147 ( .A(n4227), .B(n4161), .Z(n4397));
  AN2 U4148 ( .A(po004), .B(n4398), .Z(n4393));
  OR2 U4149 ( .A(n4399), .B(n4400), .Z(n4398));
  OR2 U4150 ( .A(n4401), .B(n4402), .Z(n4400));
  AN2 U4151 ( .A(n4310), .B(n4403), .Z(n4402));
  AN2 U4152 ( .A(n4404), .B(n4227), .Z(n4401));
  AN2 U4153 ( .A(n4405), .B(n4406), .Z(n4399));
  AN2 U4154 ( .A(n4407), .B(n3261), .Z(n4405));
  OR2 U4155 ( .A(n4408), .B(n4409), .Z(n4407));
  AN2 U4156 ( .A(n4028), .B(pi065), .Z(n4409));
  AN2 U4157 ( .A(po040), .B(n4410), .Z(n4408));
  OR2 U4158 ( .A(n4411), .B(n4412), .Z(n4410));
  AN2 U4159 ( .A(pi065), .B(n4045), .Z(n4412));
  AN2 U4160 ( .A(n4046), .B(n4156), .Z(n4411));
  OR2 U4161 ( .A(n4413), .B(n4414), .Z(po046));
  OR2 U4162 ( .A(n4415), .B(n4416), .Z(n4414));
  AN2 U4163 ( .A(n3339), .B(n4417), .Z(n4416));
  AN2 U4164 ( .A(n3341), .B(n4418), .Z(n4415));
  OR2 U4165 ( .A(n4419), .B(n4420), .Z(n4413));
  AN2 U4166 ( .A(n4421), .B(pi192), .Z(n4420));
  OR2 U4167 ( .A(n4422), .B(n4423), .Z(n4421));
  AN2 U4168 ( .A(n4424), .B(pi098), .Z(n4423));
  AN2 U4169 ( .A(n4425), .B(n4426), .Z(n4424));
  OR2 U4170 ( .A(n3242), .B(n3657), .Z(n4425));
  IV2 U4171 ( .A(n3635), .Z(n3657));
  AN2 U4172 ( .A(n4427), .B(n3638), .Z(n4422));
  OR2 U4173 ( .A(n4428), .B(n4429), .Z(n4427));
  AN2 U4174 ( .A(n4430), .B(pi171), .Z(n4429));
  AN2 U4175 ( .A(n4431), .B(n4001), .Z(n4428));
  AN2 U4176 ( .A(n4432), .B(n2837), .Z(n4419));
  OR2 U4177 ( .A(n4433), .B(n4434), .Z(n4432));
  AN2 U4178 ( .A(n4435), .B(pi003), .Z(n4434));
  AN2 U4179 ( .A(n4436), .B(n4426), .Z(n4435));
  OR2 U4180 ( .A(n3244), .B(n3616), .Z(n4436));
  IV2 U4181 ( .A(n3593), .Z(n3616));
  AN2 U4182 ( .A(n4437), .B(n3597), .Z(n4433));
  OR2 U4183 ( .A(n4438), .B(n4439), .Z(n4437));
  AN2 U4184 ( .A(n4430), .B(pi142), .Z(n4439));
  AN2 U4185 ( .A(n4431), .B(n4440), .Z(n4438));
  AN2 U4186 ( .A(n3236), .B(n4441), .Z(n4431));
  OR2 U4187 ( .A(n4442), .B(n4443), .Z(po045));
  AN2 U4188 ( .A(n4444), .B(n4445), .Z(n4443));
  OR2 U4189 ( .A(n4446), .B(n3756), .Z(n4445));
  AN2 U4190 ( .A(n4006), .B(n4005), .Z(n4446));
  OR2 U4191 ( .A(n4447), .B(n4448), .Z(n4005));
  AN2 U4192 ( .A(n4449), .B(n3301), .Z(n4447));
  AN2 U4193 ( .A(n4450), .B(n3306), .Z(n4449));
  AN2 U4194 ( .A(n3757), .B(n4451), .Z(n4442));
  OR2 U4195 ( .A(n4452), .B(n4453), .Z(n4451));
  OR2 U4196 ( .A(n4454), .B(n4455), .Z(n4453));
  AN2 U4197 ( .A(po092), .B(n4456), .Z(n4455));
  OR2 U4198 ( .A(n4008), .B(n4004), .Z(n4456));
  AN2 U4199 ( .A(n4457), .B(n4458), .Z(n4008));
  AN2 U4200 ( .A(n4458), .B(n4459), .Z(n4454));
  OR2 U4201 ( .A(n4460), .B(n4461), .Z(n4459));
  AN2 U4202 ( .A(n4462), .B(n4463), .Z(n4461));
  AN2 U4203 ( .A(n4464), .B(n4465), .Z(n4462));
  AN2 U4204 ( .A(n4466), .B(n4467), .Z(n4460));
  AN2 U4205 ( .A(n4468), .B(n4469), .Z(n4466));
  OR2 U4206 ( .A(n4470), .B(n4471), .Z(po043));
  OR2 U4207 ( .A(n4472), .B(n4473), .Z(n4471));
  AN2 U4208 ( .A(n4474), .B(n4475), .Z(n4473));
  AN2 U4209 ( .A(n4476), .B(n4337), .Z(n4474));
  AN2 U4210 ( .A(n4477), .B(n4478), .Z(n4472));
  OR2 U4211 ( .A(n4479), .B(n4480), .Z(n4477));
  AN2 U4212 ( .A(n4337), .B(n4481), .Z(n4480));
  IV2 U4213 ( .A(n4342), .Z(n4337));
  AN2 U4214 ( .A(n4342), .B(n4476), .Z(n4479));
  IV2 U4215 ( .A(n4481), .Z(n4476));
  AN2 U4216 ( .A(n4482), .B(n4481), .Z(n4470));
  OR2 U4217 ( .A(n4483), .B(n4484), .Z(n4481));
  OR2 U4218 ( .A(n4485), .B(n4486), .Z(n4484));
  AN2 U4219 ( .A(n4487), .B(n4078), .Z(n4486));
  OR2 U4220 ( .A(n4488), .B(n4489), .Z(n4487));
  AN2 U4221 ( .A(n4490), .B(n3778), .Z(n4489));
  AN2 U4222 ( .A(n3773), .B(n4491), .Z(n4488));
  AN2 U4223 ( .A(n4492), .B(n4066), .Z(n4485));
  AN2 U4224 ( .A(n4490), .B(n3773), .Z(n4492));
  AN2 U4225 ( .A(n4491), .B(n4341), .Z(n4483));
  IV2 U4226 ( .A(n4490), .Z(n4491));
  OR2 U4227 ( .A(n4493), .B(n4494), .Z(n4490));
  IV2 U4228 ( .A(n4495), .Z(n4494));
  OR2 U4229 ( .A(n4496), .B(n4497), .Z(n4495));
  AN2 U4230 ( .A(n4497), .B(n4496), .Z(n4493));
  AN2 U4231 ( .A(n4498), .B(n4499), .Z(n4496));
  IV2 U4232 ( .A(n4500), .Z(n4499));
  AN2 U4233 ( .A(n4333), .B(n4501), .Z(n4500));
  OR2 U4234 ( .A(n4501), .B(n4333), .Z(n4498));
  OR2 U4235 ( .A(n4502), .B(n4503), .Z(n4501));
  OR2 U4236 ( .A(n4504), .B(n4505), .Z(n4503));
  OR2 U4237 ( .A(n4506), .B(n4507), .Z(n4505));
  AN2 U4238 ( .A(n4508), .B(n4509), .Z(n4507));
  AN2 U4239 ( .A(n4510), .B(n4511), .Z(n4506));
  AN2 U4240 ( .A(n4512), .B(n4513), .Z(n4504));
  OR2 U4241 ( .A(n4514), .B(n4515), .Z(n4502));
  AN2 U4242 ( .A(n4516), .B(n4517), .Z(n4515));
  AN2 U4243 ( .A(po102), .B(n4518), .Z(n4514));
  OR2 U4244 ( .A(n4519), .B(n4520), .Z(n4518));
  AN2 U4245 ( .A(n4513), .B(n4521), .Z(n4520));
  OR2 U4246 ( .A(n4522), .B(n4523), .Z(n4513));
  AN2 U4247 ( .A(n4508), .B(n3773), .Z(n4523));
  AN2 U4248 ( .A(po025), .B(n4516), .Z(n4522));
  AN2 U4249 ( .A(n4508), .B(n4524), .Z(n4519));
  IV2 U4250 ( .A(n4510), .Z(n4508));
  OR2 U4251 ( .A(n4525), .B(n4526), .Z(n4510));
  AN2 U4252 ( .A(n4527), .B(n4528), .Z(n4526));
  OR2 U4253 ( .A(n4529), .B(n4530), .Z(n4527));
  OR2 U4254 ( .A(n4531), .B(n4532), .Z(n4530));
  AN2 U4255 ( .A(po025), .B(n4533), .Z(n4532));
  OR2 U4256 ( .A(n4534), .B(n4535), .Z(n4533));
  OR2 U4257 ( .A(n4356), .B(n4536), .Z(n4535));
  AN2 U4258 ( .A(n4537), .B(n4538), .Z(n4536));
  AN2 U4259 ( .A(n4539), .B(n4540), .Z(n4537));
  AN2 U4260 ( .A(n3890), .B(n4541), .Z(n4534));
  OR2 U4261 ( .A(n4542), .B(n4543), .Z(n4541));
  AN2 U4262 ( .A(n4085), .B(n4544), .Z(n4542));
  AN2 U4263 ( .A(n3778), .B(n4545), .Z(n4531));
  OR2 U4264 ( .A(n4546), .B(n4547), .Z(n4545));
  OR2 U4265 ( .A(n4548), .B(n4549), .Z(n4547));
  AN2 U4266 ( .A(n3775), .B(n4550), .Z(n4549));
  AN2 U4267 ( .A(n4524), .B(n4333), .Z(n4548));
  AN2 U4268 ( .A(n4086), .B(n4551), .Z(n4546));
  OR2 U4269 ( .A(n4552), .B(n4553), .Z(n4529));
  AN2 U4270 ( .A(n4554), .B(n4555), .Z(n4553));
  OR2 U4271 ( .A(n4556), .B(n3888), .Z(n4555));
  AN2 U4272 ( .A(pi192), .B(n4557), .Z(n4556));
  AN2 U4273 ( .A(n4558), .B(n4559), .Z(n4554));
  OR2 U4274 ( .A(n4085), .B(n4560), .Z(n4558));
  AN2 U4275 ( .A(n4561), .B(n3773), .Z(n4560));
  AN2 U4276 ( .A(n4562), .B(n4563), .Z(n4552));
  OR2 U4277 ( .A(n4564), .B(n4565), .Z(n4563));
  AN2 U4278 ( .A(n4566), .B(n4567), .Z(n4564));
  AN2 U4279 ( .A(n3773), .B(n4076), .Z(n4566));
  OR2 U4280 ( .A(pi076), .B(n4557), .Z(n4562));
  AN2 U4281 ( .A(n4516), .B(n4568), .Z(n4525));
  OR2 U4282 ( .A(n4569), .B(n4570), .Z(n4568));
  OR2 U4283 ( .A(n4571), .B(n4572), .Z(n4570));
  OR2 U4284 ( .A(n4573), .B(n4574), .Z(n4572));
  AN2 U4285 ( .A(n4575), .B(n4576), .Z(n4574));
  AN2 U4286 ( .A(n4577), .B(n4076), .Z(n4575));
  AN2 U4287 ( .A(n3773), .B(n4578), .Z(n4577));
  AN2 U4288 ( .A(n4579), .B(n4580), .Z(n4573));
  OR2 U4289 ( .A(n4581), .B(n4565), .Z(n4579));
  AN2 U4290 ( .A(n4539), .B(n4582), .Z(n4565));
  AN2 U4291 ( .A(n2837), .B(n4550), .Z(n4582));
  IV2 U4292 ( .A(n4540), .Z(n4550));
  AN2 U4293 ( .A(n4567), .B(n4076), .Z(n4581));
  AN2 U4294 ( .A(n4086), .B(n4583), .Z(n4571));
  OR2 U4295 ( .A(n4584), .B(n4585), .Z(n4583));
  AN2 U4296 ( .A(n4543), .B(n3773), .Z(n4585));
  AN2 U4297 ( .A(n4586), .B(n4544), .Z(n4584));
  OR2 U4298 ( .A(n4085), .B(n3778), .Z(n4586));
  AN2 U4299 ( .A(n4557), .B(n3888), .Z(n4086));
  OR2 U4300 ( .A(n4587), .B(n4588), .Z(n4569));
  AN2 U4301 ( .A(n4589), .B(n4590), .Z(n4588));
  OR2 U4302 ( .A(n4591), .B(n3890), .Z(n4590));
  AN2 U4303 ( .A(po025), .B(pi192), .Z(n4591));
  AN2 U4304 ( .A(n4559), .B(n4592), .Z(n4589));
  OR2 U4305 ( .A(n4561), .B(n4085), .Z(n4592));
  OR2 U4306 ( .A(n4551), .B(n4353), .Z(n4559));
  AN2 U4307 ( .A(n4593), .B(n3775), .Z(n4587));
  AN2 U4308 ( .A(n2837), .B(n4576), .Z(n3775));
  AN2 U4309 ( .A(n4594), .B(n4540), .Z(n4593));
  OR2 U4310 ( .A(n4567), .B(n4066), .Z(n4540));
  OR2 U4311 ( .A(n4539), .B(n3778), .Z(n4594));
  IV2 U4312 ( .A(n4528), .Z(n4516));
  OR2 U4313 ( .A(n4595), .B(n4596), .Z(n4497));
  AN2 U4314 ( .A(n4597), .B(n4598), .Z(n4596));
  OR2 U4315 ( .A(n4599), .B(n4600), .Z(n4598));
  AN2 U4316 ( .A(n4601), .B(n4602), .Z(n4600));
  IV2 U4317 ( .A(n4603), .Z(n4599));
  OR2 U4318 ( .A(n4602), .B(n4601), .Z(n4603));
  OR2 U4319 ( .A(n4604), .B(n4605), .Z(n4601));
  AN2 U4320 ( .A(n3295), .B(n4606), .Z(n4605));
  AN2 U4321 ( .A(n4450), .B(n3301), .Z(n4604));
  AN2 U4322 ( .A(n4607), .B(n4608), .Z(n4602));
  OR2 U4323 ( .A(n4609), .B(n4610), .Z(n4608));
  IV2 U4324 ( .A(n4611), .Z(n4610));
  OR2 U4325 ( .A(n4611), .B(n4612), .Z(n4607));
  IV2 U4326 ( .A(n4609), .Z(n4612));
  OR2 U4327 ( .A(n4613), .B(n4614), .Z(n4609));
  OR2 U4328 ( .A(n4615), .B(n4616), .Z(n4614));
  AN2 U4329 ( .A(n4004), .B(n4617), .Z(n4616));
  OR2 U4330 ( .A(n4618), .B(n4619), .Z(n4617));
  AN2 U4331 ( .A(n4620), .B(n4463), .Z(n4619));
  AN2 U4332 ( .A(n4621), .B(n4464), .Z(n4620));
  AN2 U4333 ( .A(n4622), .B(n4467), .Z(n4618));
  AN2 U4334 ( .A(n4623), .B(n4468), .Z(n4622));
  AN2 U4335 ( .A(n4006), .B(n4624), .Z(n4615));
  OR2 U4336 ( .A(n4625), .B(n4626), .Z(n4613));
  AN2 U4337 ( .A(n4627), .B(n4628), .Z(n4626));
  OR2 U4338 ( .A(n4629), .B(n4630), .Z(n4627));
  AN2 U4339 ( .A(n4631), .B(pi192), .Z(n4630));
  AN2 U4340 ( .A(n4632), .B(pi158), .Z(n4631));
  AN2 U4341 ( .A(n4633), .B(n4634), .Z(n4632));
  OR2 U4342 ( .A(n4635), .B(n4465), .Z(n4634));
  OR2 U4343 ( .A(n4464), .B(n4636), .Z(n4633));
  OR2 U4344 ( .A(n4621), .B(n3301), .Z(n4636));
  AN2 U4345 ( .A(n4637), .B(n2837), .Z(n4629));
  AN2 U4346 ( .A(n4638), .B(pi151), .Z(n4637));
  AN2 U4347 ( .A(n4639), .B(n4640), .Z(n4638));
  OR2 U4348 ( .A(n4641), .B(n4469), .Z(n4640));
  OR2 U4349 ( .A(n4468), .B(n4642), .Z(n4639));
  OR2 U4350 ( .A(n4623), .B(n3301), .Z(n4642));
  AN2 U4351 ( .A(n4643), .B(po092), .Z(n4625));
  AN2 U4352 ( .A(n4644), .B(n3295), .Z(n4643));
  AN2 U4353 ( .A(n4645), .B(n4646), .Z(n4644));
  OR2 U4354 ( .A(pi192), .B(n4647), .Z(n4646));
  AN2 U4355 ( .A(n4641), .B(n4648), .Z(n4647));
  OR2 U4356 ( .A(n2837), .B(n4649), .Z(n4645));
  AN2 U4357 ( .A(n4635), .B(n3908), .Z(n4649));
  IV2 U4358 ( .A(n3761), .Z(n4597));
  AN2 U4359 ( .A(n4650), .B(n3761), .Z(n4595));
  OR2 U4360 ( .A(n4651), .B(n4652), .Z(n3761));
  AN2 U4361 ( .A(n4653), .B(n4654), .Z(n4651));
  AN2 U4362 ( .A(n4333), .B(n4528), .Z(n4654));
  OR2 U4363 ( .A(n4655), .B(n4656), .Z(n4528));
  AN2 U4364 ( .A(n4657), .B(n3083), .Z(n4655));
  AN2 U4365 ( .A(n3018), .B(n4658), .Z(n4657));
  OR2 U4366 ( .A(n4659), .B(n4660), .Z(n4658));
  OR2 U4367 ( .A(n4661), .B(n4662), .Z(n4660));
  AN2 U4368 ( .A(n4663), .B(n3010), .Z(n4662));
  AN2 U4369 ( .A(n4664), .B(n3049), .Z(n4661));
  OR2 U4370 ( .A(n4665), .B(n4663), .Z(n4664));
  AN2 U4371 ( .A(n4666), .B(n3010), .Z(n4665));
  OR2 U4372 ( .A(n3100), .B(n4667), .Z(n4659));
  AN2 U4373 ( .A(n4668), .B(n3012), .Z(n4667));
  OR2 U4374 ( .A(n4669), .B(n4670), .Z(n4668));
  AN2 U4375 ( .A(n4671), .B(pi201), .Z(n4670));
  AN2 U4376 ( .A(n4672), .B(n3115), .Z(n4671));
  OR2 U4377 ( .A(n4673), .B(n3173), .Z(n4672));
  AN2 U4378 ( .A(n2837), .B(n3049), .Z(n4673));
  AN2 U4379 ( .A(n4674), .B(pi088), .Z(n4669));
  AN2 U4380 ( .A(n4675), .B(n3108), .Z(n4674));
  OR2 U4381 ( .A(n4676), .B(n3064), .Z(n4675));
  AN2 U4382 ( .A(pi192), .B(n3049), .Z(n4676));
  AN2 U4383 ( .A(n4341), .B(n4482), .Z(n4653));
  OR2 U4384 ( .A(n4677), .B(n4678), .Z(n4650));
  OR2 U4385 ( .A(n4679), .B(n4680), .Z(n4678));
  OR2 U4386 ( .A(n4681), .B(n4682), .Z(n4680));
  AN2 U4387 ( .A(n4683), .B(n4684), .Z(n4682));
  AN2 U4388 ( .A(n4685), .B(n4648), .Z(n4683));
  AN2 U4389 ( .A(n4686), .B(n4687), .Z(n4681));
  OR2 U4390 ( .A(n4688), .B(n4689), .Z(n4687));
  OR2 U4391 ( .A(n4690), .B(n4691), .Z(n4689));
  AN2 U4392 ( .A(n4692), .B(n4621), .Z(n4691));
  AN2 U4393 ( .A(n4685), .B(n4623), .Z(n4690));
  AN2 U4394 ( .A(n4693), .B(n3300), .Z(n4688));
  IV2 U4395 ( .A(n4684), .Z(n4686));
  OR2 U4396 ( .A(n4694), .B(n4695), .Z(n4679));
  AN2 U4397 ( .A(n4696), .B(n3300), .Z(n4695));
  AN2 U4398 ( .A(po014), .B(n4684), .Z(n4696));
  OR2 U4399 ( .A(n4697), .B(n4698), .Z(n4684));
  AN2 U4400 ( .A(n4699), .B(n4450), .Z(n4697));
  AN2 U4401 ( .A(po039), .B(n4700), .Z(n4694));
  OR2 U4402 ( .A(n4701), .B(n4702), .Z(n4700));
  AN2 U4403 ( .A(n4698), .B(n4703), .Z(n4702));
  AN2 U4404 ( .A(n4704), .B(n4606), .Z(n4698));
  AN2 U4405 ( .A(n4705), .B(n4706), .Z(n4701));
  AN2 U4406 ( .A(n4707), .B(n4708), .Z(n4705));
  OR2 U4407 ( .A(n4704), .B(n3295), .Z(n4708));
  OR2 U4408 ( .A(n4699), .B(n3301), .Z(n4707));
  OR2 U4409 ( .A(n4709), .B(n4710), .Z(n4677));
  AN2 U4410 ( .A(n4711), .B(n4699), .Z(n4710));
  IV2 U4411 ( .A(n4704), .Z(n4699));
  AN2 U4412 ( .A(n4450), .B(n4712), .Z(n4711));
  OR2 U4413 ( .A(po014), .B(n3301), .Z(n4712));
  AN2 U4414 ( .A(n4713), .B(n4704), .Z(n4709));
  OR2 U4415 ( .A(n4714), .B(n4715), .Z(n4704));
  OR2 U4416 ( .A(n4716), .B(n4717), .Z(n4715));
  OR2 U4417 ( .A(n4718), .B(n4719), .Z(n4717));
  IV2 U4418 ( .A(n4720), .Z(n4719));
  OR2 U4419 ( .A(n4721), .B(n4006), .Z(n4720));
  OR2 U4420 ( .A(n4444), .B(n3756), .Z(n4721));
  AN2 U4421 ( .A(n4722), .B(n4006), .Z(n4718));
  AN2 U4422 ( .A(n4444), .B(n4452), .Z(n4722));
  OR2 U4423 ( .A(n4723), .B(n4724), .Z(n4452));
  OR2 U4424 ( .A(n4725), .B(n4726), .Z(n4724));
  AN2 U4425 ( .A(po092), .B(n4009), .Z(n4726));
  OR2 U4426 ( .A(n4727), .B(n4728), .Z(n4009));
  AN2 U4427 ( .A(n3295), .B(n4729), .Z(n4728));
  AN2 U4428 ( .A(n4606), .B(n4457), .Z(n4727));
  OR2 U4429 ( .A(n4730), .B(n4706), .Z(n4457));
  OR2 U4430 ( .A(n4731), .B(n4732), .Z(n4706));
  AN2 U4431 ( .A(n4733), .B(pi192), .Z(n4732));
  AN2 U4432 ( .A(n4465), .B(n3870), .Z(n4733));
  AN2 U4433 ( .A(n4734), .B(n2837), .Z(n4731));
  AN2 U4434 ( .A(n4469), .B(n4735), .Z(n4734));
  AN2 U4435 ( .A(po039), .B(n4729), .Z(n4730));
  OR2 U4436 ( .A(po014), .B(n4736), .Z(n4729));
  AN2 U4437 ( .A(n4737), .B(n4606), .Z(n4725));
  AN2 U4438 ( .A(po014), .B(n4738), .Z(n4737));
  OR2 U4439 ( .A(n4739), .B(n4740), .Z(n4738));
  AN2 U4440 ( .A(n4463), .B(n4464), .Z(n4740));
  AN2 U4441 ( .A(n4467), .B(n4468), .Z(n4739));
  OR2 U4442 ( .A(n4741), .B(n4742), .Z(n4723));
  AN2 U4443 ( .A(n4743), .B(n4463), .Z(n4742));
  AN2 U4444 ( .A(n3909), .B(pi192), .Z(n4463));
  IV2 U4445 ( .A(pi158), .Z(n3909));
  AN2 U4446 ( .A(n4744), .B(n3908), .Z(n4743));
  OR2 U4447 ( .A(n4745), .B(n3295), .Z(n4744));
  AN2 U4448 ( .A(n4606), .B(n4464), .Z(n4745));
  AN2 U4449 ( .A(n4746), .B(n4467), .Z(n4741));
  AN2 U4450 ( .A(n2837), .B(n4747), .Z(n4467));
  AN2 U4451 ( .A(n4748), .B(n4648), .Z(n4746));
  OR2 U4452 ( .A(n4749), .B(n3295), .Z(n4748));
  AN2 U4453 ( .A(n4606), .B(n4468), .Z(n4749));
  AN2 U4454 ( .A(n3756), .B(n4611), .Z(n4716));
  OR2 U4455 ( .A(n4750), .B(n4751), .Z(n4611));
  AN2 U4456 ( .A(n4004), .B(n4444), .Z(n4750));
  IV2 U4457 ( .A(n4006), .Z(n4004));
  AN2 U4458 ( .A(n4628), .B(n4752), .Z(n3756));
  OR2 U4459 ( .A(n3758), .B(n3760), .Z(n4714));
  AN2 U4460 ( .A(n4448), .B(n4751), .Z(n3758));
  OR2 U4461 ( .A(n4713), .B(n4693), .Z(n4448));
  OR2 U4462 ( .A(n4753), .B(n4754), .Z(n4693));
  AN2 U4463 ( .A(n4621), .B(pi192), .Z(n4754));
  AN2 U4464 ( .A(n4623), .B(n2837), .Z(n4753));
  AN2 U4465 ( .A(n3301), .B(n4624), .Z(n4713));
  OR2 U4466 ( .A(n4755), .B(n4756), .Z(po042));
  AN2 U4467 ( .A(n4757), .B(n2837), .Z(n4756));
  OR2 U4468 ( .A(n4758), .B(n4759), .Z(n4757));
  OR2 U4469 ( .A(n4760), .B(n4761), .Z(n4759));
  AN2 U4470 ( .A(n4762), .B(n4763), .Z(n4761));
  OR2 U4471 ( .A(n4764), .B(n4765), .Z(n4763));
  IV2 U4472 ( .A(n4766), .Z(n4762));
  AN2 U4473 ( .A(n4765), .B(n4764), .Z(n4766));
  OR2 U4474 ( .A(n4767), .B(n4768), .Z(n4764));
  AN2 U4475 ( .A(n4769), .B(n4770), .Z(n4768));
  AN2 U4476 ( .A(n4771), .B(pi028), .Z(n4767));
  AN2 U4477 ( .A(n4772), .B(n4773), .Z(n4765));
  OR2 U4478 ( .A(n4774), .B(pi094), .Z(n4773));
  IV2 U4479 ( .A(n4775), .Z(n4772));
  AN2 U4480 ( .A(n4774), .B(pi094), .Z(n4775));
  AN2 U4481 ( .A(n4776), .B(n4777), .Z(n4774));
  OR2 U4482 ( .A(n4778), .B(pi173), .Z(n4777));
  OR2 U4483 ( .A(n4779), .B(pi163), .Z(n4776));
  IV2 U4484 ( .A(pi173), .Z(n4779));
  AN2 U4485 ( .A(n4780), .B(n4781), .Z(n4760));
  IV2 U4486 ( .A(n4782), .Z(n4781));
  AN2 U4487 ( .A(n4783), .B(n4784), .Z(n4782));
  OR2 U4488 ( .A(n4784), .B(n4783), .Z(n4780));
  AN2 U4489 ( .A(n4785), .B(n4786), .Z(n4783));
  IV2 U4490 ( .A(n4787), .Z(n4786));
  AN2 U4491 ( .A(n4788), .B(n4789), .Z(n4787));
  OR2 U4492 ( .A(n4789), .B(n4788), .Z(n4785));
  OR2 U4493 ( .A(n4790), .B(n4791), .Z(n4788));
  AN2 U4494 ( .A(pi025), .B(n4792), .Z(n4791));
  IV2 U4495 ( .A(n4793), .Z(n4790));
  OR2 U4496 ( .A(n4792), .B(pi025), .Z(n4793));
  IV2 U4497 ( .A(pi035), .Z(n4792));
  AN2 U4498 ( .A(n4794), .B(n4795), .Z(n4789));
  IV2 U4499 ( .A(n4796), .Z(n4795));
  AN2 U4500 ( .A(pi056), .B(n4797), .Z(n4796));
  OR2 U4501 ( .A(n4797), .B(pi056), .Z(n4794));
  IV2 U4502 ( .A(pi100), .Z(n4797));
  OR2 U4503 ( .A(n4798), .B(n4799), .Z(n4784));
  IV2 U4504 ( .A(n4800), .Z(n4799));
  OR2 U4505 ( .A(n4801), .B(n4802), .Z(n4800));
  AN2 U4506 ( .A(n4802), .B(n4801), .Z(n4798));
  AN2 U4507 ( .A(n4803), .B(n4804), .Z(n4801));
  IV2 U4508 ( .A(n4805), .Z(n4804));
  AN2 U4509 ( .A(pi126), .B(n4806), .Z(n4805));
  OR2 U4510 ( .A(n4806), .B(pi126), .Z(n4803));
  IV2 U4511 ( .A(pi146), .Z(n4806));
  OR2 U4512 ( .A(n4807), .B(n4808), .Z(n4802));
  AN2 U4513 ( .A(pi190), .B(n4809), .Z(n4808));
  IV2 U4514 ( .A(pi202), .Z(n4809));
  AN2 U4515 ( .A(pi202), .B(n4810), .Z(n4807));
  IV2 U4516 ( .A(pi190), .Z(n4810));
  OR2 U4517 ( .A(n4811), .B(n4812), .Z(n4758));
  AN2 U4518 ( .A(n4813), .B(n4814), .Z(n4812));
  IV2 U4519 ( .A(n4815), .Z(n4814));
  AN2 U4520 ( .A(n4816), .B(n4817), .Z(n4815));
  OR2 U4521 ( .A(n4817), .B(n4816), .Z(n4813));
  AN2 U4522 ( .A(n4818), .B(n4819), .Z(n4816));
  OR2 U4523 ( .A(n4820), .B(pi019), .Z(n4819));
  OR2 U4524 ( .A(n4821), .B(n4822), .Z(n4818));
  IV2 U4525 ( .A(pi019), .Z(n4822));
  OR2 U4526 ( .A(n4823), .B(n4824), .Z(n4817));
  IV2 U4527 ( .A(n4825), .Z(n4824));
  OR2 U4528 ( .A(n4826), .B(pi085), .Z(n4825));
  AN2 U4529 ( .A(n4826), .B(pi085), .Z(n4823));
  AN2 U4530 ( .A(n4827), .B(n4828), .Z(n4826));
  OR2 U4531 ( .A(n4829), .B(pi167), .Z(n4828));
  IV2 U4532 ( .A(pi110), .Z(n4829));
  OR2 U4533 ( .A(n4830), .B(pi110), .Z(n4827));
  IV2 U4534 ( .A(pi167), .Z(n4830));
  AN2 U4535 ( .A(n4831), .B(n4832), .Z(n4811));
  IV2 U4536 ( .A(n4833), .Z(n4832));
  AN2 U4537 ( .A(n4834), .B(n4835), .Z(n4833));
  OR2 U4538 ( .A(n4835), .B(n4834), .Z(n4831));
  AN2 U4539 ( .A(n4836), .B(n4837), .Z(n4834));
  OR2 U4540 ( .A(n4838), .B(pi020), .Z(n4837));
  OR2 U4541 ( .A(n4839), .B(n4840), .Z(n4836));
  IV2 U4542 ( .A(pi020), .Z(n4840));
  OR2 U4543 ( .A(n4841), .B(n4842), .Z(n4835));
  IV2 U4544 ( .A(n4843), .Z(n4842));
  OR2 U4545 ( .A(n4844), .B(pi047), .Z(n4843));
  AN2 U4546 ( .A(n4844), .B(pi047), .Z(n4841));
  AN2 U4547 ( .A(n4845), .B(n4846), .Z(n4844));
  OR2 U4548 ( .A(n4847), .B(pi153), .Z(n4846));
  IV2 U4549 ( .A(pi075), .Z(n4847));
  OR2 U4550 ( .A(n4848), .B(pi075), .Z(n4845));
  IV2 U4551 ( .A(pi153), .Z(n4848));
  AN2 U4552 ( .A(pi192), .B(n4849), .Z(n4755));
  OR2 U4553 ( .A(n4850), .B(n4851), .Z(n4849));
  OR2 U4554 ( .A(n4852), .B(n4853), .Z(n4851));
  AN2 U4555 ( .A(n4854), .B(n4855), .Z(n4853));
  OR2 U4556 ( .A(n4856), .B(n4857), .Z(n4855));
  IV2 U4557 ( .A(n4858), .Z(n4854));
  AN2 U4558 ( .A(n4857), .B(n4856), .Z(n4858));
  OR2 U4559 ( .A(n4859), .B(n4860), .Z(n4856));
  AN2 U4560 ( .A(n4839), .B(n4861), .Z(n4860));
  AN2 U4561 ( .A(n4838), .B(po014), .Z(n4859));
  IV2 U4562 ( .A(n4839), .Z(n4838));
  OR2 U4563 ( .A(n4862), .B(n4863), .Z(n4839));
  AN2 U4564 ( .A(n4864), .B(pi192), .Z(n4863));
  OR2 U4565 ( .A(n4865), .B(n4866), .Z(n4864));
  IV2 U4566 ( .A(n4867), .Z(n4866));
  OR2 U4567 ( .A(n4868), .B(n4869), .Z(n4867));
  AN2 U4568 ( .A(n4869), .B(n4868), .Z(n4865));
  AN2 U4569 ( .A(n4870), .B(n4871), .Z(n4868));
  OR2 U4570 ( .A(n4872), .B(po024), .Z(n4871));
  IV2 U4571 ( .A(n4873), .Z(n4872));
  OR2 U4572 ( .A(n4873), .B(n4874), .Z(n4870));
  OR2 U4573 ( .A(n4875), .B(n4876), .Z(n4873));
  AN2 U4574 ( .A(po025), .B(n4877), .Z(n4876));
  AN2 U4575 ( .A(po059), .B(n4557), .Z(n4875));
  OR2 U4576 ( .A(n4878), .B(n4879), .Z(n4869));
  AN2 U4577 ( .A(n4880), .B(n4881), .Z(n4879));
  AN2 U4578 ( .A(n4882), .B(po072), .Z(n4878));
  IV2 U4579 ( .A(n4880), .Z(n4882));
  OR2 U4580 ( .A(n4883), .B(n4884), .Z(n4880));
  AN2 U4581 ( .A(po084), .B(n4885), .Z(n4884));
  AN2 U4582 ( .A(po102), .B(n4886), .Z(n4883));
  IV2 U4583 ( .A(po084), .Z(n4886));
  AN2 U4584 ( .A(n4887), .B(n2837), .Z(n4862));
  OR2 U4585 ( .A(n4888), .B(n4889), .Z(n4887));
  AN2 U4586 ( .A(n4890), .B(n4891), .Z(n4889));
  IV2 U4587 ( .A(n4892), .Z(n4888));
  OR2 U4588 ( .A(n4891), .B(n4890), .Z(n4892));
  OR2 U4589 ( .A(n4893), .B(n4894), .Z(n4890));
  IV2 U4590 ( .A(n4895), .Z(n4894));
  OR2 U4591 ( .A(n4896), .B(pi014), .Z(n4895));
  AN2 U4592 ( .A(n4896), .B(pi014), .Z(n4893));
  AN2 U4593 ( .A(n4897), .B(n4898), .Z(n4896));
  OR2 U4594 ( .A(n4899), .B(pi111), .Z(n4898));
  OR2 U4595 ( .A(n4900), .B(pi097), .Z(n4897));
  IV2 U4596 ( .A(pi111), .Z(n4900));
  AN2 U4597 ( .A(n4901), .B(n4902), .Z(n4891));
  OR2 U4598 ( .A(n4903), .B(pi143), .Z(n4902));
  IV2 U4599 ( .A(n4904), .Z(n4901));
  AN2 U4600 ( .A(n4903), .B(pi143), .Z(n4904));
  AN2 U4601 ( .A(n4905), .B(n4906), .Z(n4903));
  OR2 U4602 ( .A(n4907), .B(pi189), .Z(n4906));
  IV2 U4603 ( .A(n4908), .Z(n4905));
  AN2 U4604 ( .A(pi189), .B(n4907), .Z(n4908));
  IV2 U4605 ( .A(pi176), .Z(n4907));
  AN2 U4606 ( .A(n4909), .B(n4910), .Z(n4857));
  OR2 U4607 ( .A(n4911), .B(po039), .Z(n4910));
  IV2 U4608 ( .A(n4912), .Z(n4911));
  OR2 U4609 ( .A(n4912), .B(n3300), .Z(n4909));
  OR2 U4610 ( .A(n4913), .B(n4914), .Z(n4912));
  AN2 U4611 ( .A(po063), .B(n4628), .Z(n4914));
  AN2 U4612 ( .A(po092), .B(n4915), .Z(n4913));
  AN2 U4613 ( .A(n4916), .B(n4917), .Z(n4852));
  IV2 U4614 ( .A(n4918), .Z(n4917));
  AN2 U4615 ( .A(n4919), .B(n4920), .Z(n4918));
  OR2 U4616 ( .A(n4920), .B(n4919), .Z(n4916));
  IV2 U4617 ( .A(n4921), .Z(n4919));
  OR2 U4618 ( .A(n4922), .B(n4923), .Z(n4921));
  AN2 U4619 ( .A(n4821), .B(n3391), .Z(n4923));
  IV2 U4620 ( .A(n4924), .Z(n3391));
  AN2 U4621 ( .A(n4924), .B(n4820), .Z(n4922));
  IV2 U4622 ( .A(n4821), .Z(n4820));
  OR2 U4623 ( .A(n4925), .B(n4926), .Z(n4821));
  AN2 U4624 ( .A(n4927), .B(pi192), .Z(n4926));
  OR2 U4625 ( .A(n4928), .B(n4929), .Z(n4927));
  IV2 U4626 ( .A(n4930), .Z(n4929));
  OR2 U4627 ( .A(n4931), .B(n4932), .Z(n4930));
  AN2 U4628 ( .A(n4932), .B(n4931), .Z(n4928));
  AN2 U4629 ( .A(n4933), .B(n4934), .Z(n4931));
  OR2 U4630 ( .A(n4935), .B(po001), .Z(n4934));
  IV2 U4631 ( .A(n4936), .Z(n4935));
  OR2 U4632 ( .A(n4936), .B(n4937), .Z(n4933));
  OR2 U4633 ( .A(n4938), .B(n4939), .Z(n4936));
  AN2 U4634 ( .A(po011), .B(n4441), .Z(n4939));
  AN2 U4635 ( .A(po036), .B(n3688), .Z(n4938));
  OR2 U4636 ( .A(n4940), .B(n4941), .Z(n4932));
  AN2 U4637 ( .A(n4942), .B(n4943), .Z(n4941));
  AN2 U4638 ( .A(n4944), .B(po057), .Z(n4940));
  IV2 U4639 ( .A(n4942), .Z(n4944));
  OR2 U4640 ( .A(n4945), .B(n4946), .Z(n4942));
  AN2 U4641 ( .A(po069), .B(n4947), .Z(n4946));
  AN2 U4642 ( .A(po082), .B(n4948), .Z(n4945));
  IV2 U4643 ( .A(po069), .Z(n4948));
  AN2 U4644 ( .A(n4949), .B(n2837), .Z(n4925));
  OR2 U4645 ( .A(n4950), .B(n4951), .Z(n4949));
  AN2 U4646 ( .A(n4952), .B(n4953), .Z(n4951));
  IV2 U4647 ( .A(n4954), .Z(n4950));
  OR2 U4648 ( .A(n4953), .B(n4952), .Z(n4954));
  OR2 U4649 ( .A(n4955), .B(n4956), .Z(n4952));
  IV2 U4650 ( .A(n4957), .Z(n4956));
  OR2 U4651 ( .A(n4958), .B(pi024), .Z(n4957));
  AN2 U4652 ( .A(n4958), .B(pi024), .Z(n4955));
  AN2 U4653 ( .A(n4959), .B(n4960), .Z(n4958));
  OR2 U4654 ( .A(n4961), .B(pi078), .Z(n4960));
  OR2 U4655 ( .A(n4962), .B(pi030), .Z(n4959));
  IV2 U4656 ( .A(pi078), .Z(n4962));
  AN2 U4657 ( .A(n4963), .B(n4964), .Z(n4953));
  OR2 U4658 ( .A(n4965), .B(pi087), .Z(n4964));
  IV2 U4659 ( .A(n4966), .Z(n4963));
  AN2 U4660 ( .A(n4965), .B(pi087), .Z(n4966));
  AN2 U4661 ( .A(n4967), .B(n4968), .Z(n4965));
  OR2 U4662 ( .A(n4969), .B(pi164), .Z(n4968));
  OR2 U4663 ( .A(n4970), .B(pi159), .Z(n4967));
  IV2 U4664 ( .A(pi164), .Z(n4970));
  OR2 U4665 ( .A(n4971), .B(n4972), .Z(n4924));
  AN2 U4666 ( .A(po027), .B(n3512), .Z(n4972));
  AN2 U4667 ( .A(po104), .B(n3363), .Z(n4971));
  OR2 U4668 ( .A(n4973), .B(n4974), .Z(n4920));
  AN2 U4669 ( .A(po038), .B(n3380), .Z(n4974));
  AN2 U4670 ( .A(po071), .B(n4975), .Z(n4973));
  OR2 U4671 ( .A(n4976), .B(n4977), .Z(n4850));
  AN2 U4672 ( .A(n4978), .B(n4979), .Z(n4977));
  OR2 U4673 ( .A(n4980), .B(n4981), .Z(n4979));
  IV2 U4674 ( .A(n4982), .Z(n4978));
  AN2 U4675 ( .A(n4981), .B(n4980), .Z(n4982));
  OR2 U4676 ( .A(n4983), .B(n4984), .Z(n4980));
  AN2 U4677 ( .A(n4769), .B(n3049), .Z(n4984));
  AN2 U4678 ( .A(n4771), .B(po010), .Z(n4983));
  IV2 U4679 ( .A(n4769), .Z(n4771));
  OR2 U4680 ( .A(n4985), .B(n4986), .Z(n4769));
  AN2 U4681 ( .A(n4987), .B(pi192), .Z(n4986));
  OR2 U4682 ( .A(n4988), .B(n4989), .Z(n4987));
  IV2 U4683 ( .A(n4990), .Z(n4989));
  OR2 U4684 ( .A(n4991), .B(n4992), .Z(n4990));
  AN2 U4685 ( .A(n4992), .B(n4991), .Z(n4988));
  AN2 U4686 ( .A(n4993), .B(n4994), .Z(n4991));
  OR2 U4687 ( .A(n4995), .B(po031), .Z(n4994));
  IV2 U4688 ( .A(n4996), .Z(n4995));
  OR2 U4689 ( .A(n4996), .B(n2962), .Z(n4993));
  OR2 U4690 ( .A(n4997), .B(n4998), .Z(n4996));
  AN2 U4691 ( .A(po044), .B(n4999), .Z(n4998));
  IV2 U4692 ( .A(po052), .Z(n4999));
  AN2 U4693 ( .A(po052), .B(n5000), .Z(n4997));
  OR2 U4694 ( .A(n5001), .B(n5002), .Z(n4992));
  AN2 U4695 ( .A(n5003), .B(n5004), .Z(n5002));
  AN2 U4696 ( .A(n5005), .B(po079), .Z(n5001));
  IV2 U4697 ( .A(n5003), .Z(n5005));
  OR2 U4698 ( .A(n5006), .B(n5007), .Z(n5003));
  AN2 U4699 ( .A(po106), .B(n2931), .Z(n5007));
  AN2 U4700 ( .A(po107), .B(n5008), .Z(n5006));
  AN2 U4701 ( .A(n5009), .B(n2837), .Z(n4985));
  OR2 U4702 ( .A(n5010), .B(n5011), .Z(n5009));
  IV2 U4703 ( .A(n5012), .Z(n5011));
  OR2 U4704 ( .A(n5013), .B(n5014), .Z(n5012));
  AN2 U4705 ( .A(n5014), .B(n5013), .Z(n5010));
  AN2 U4706 ( .A(n5015), .B(n5016), .Z(n5013));
  OR2 U4707 ( .A(n5017), .B(pi011), .Z(n5016));
  IV2 U4708 ( .A(n5018), .Z(n5017));
  OR2 U4709 ( .A(n5018), .B(n5019), .Z(n5015));
  OR2 U4710 ( .A(n5020), .B(n5021), .Z(n5018));
  AN2 U4711 ( .A(pi021), .B(n5022), .Z(n5021));
  AN2 U4712 ( .A(pi032), .B(n5023), .Z(n5020));
  IV2 U4713 ( .A(pi021), .Z(n5023));
  OR2 U4714 ( .A(n5024), .B(n5025), .Z(n5014));
  AN2 U4715 ( .A(n5026), .B(n5027), .Z(n5025));
  AN2 U4716 ( .A(n5028), .B(pi086), .Z(n5024));
  IV2 U4717 ( .A(n5026), .Z(n5028));
  OR2 U4718 ( .A(n5029), .B(n5030), .Z(n5026));
  AN2 U4719 ( .A(pi115), .B(n5031), .Z(n5030));
  AN2 U4720 ( .A(pi165), .B(n5032), .Z(n5029));
  IV2 U4721 ( .A(pi115), .Z(n5032));
  AN2 U4722 ( .A(n5033), .B(n5034), .Z(n4981));
  OR2 U4723 ( .A(n5035), .B(po035), .Z(n5034));
  IV2 U4724 ( .A(n5036), .Z(n5035));
  OR2 U4725 ( .A(n5036), .B(n5037), .Z(n5033));
  OR2 U4726 ( .A(n5038), .B(n5039), .Z(n5036));
  AN2 U4727 ( .A(po070), .B(n3286), .Z(n5039));
  AN2 U4728 ( .A(po099), .B(n5040), .Z(n5038));
  AN2 U4729 ( .A(n5041), .B(n5042), .Z(n4976));
  OR2 U4730 ( .A(n5043), .B(n5044), .Z(n5042));
  IV2 U4731 ( .A(n5045), .Z(n5041));
  AN2 U4732 ( .A(n5044), .B(n5043), .Z(n5045));
  OR2 U4733 ( .A(n5046), .B(n5047), .Z(n5043));
  IV2 U4734 ( .A(n5048), .Z(n5047));
  OR2 U4735 ( .A(n5049), .B(n5050), .Z(n5048));
  AN2 U4736 ( .A(n5050), .B(n5049), .Z(n5046));
  AN2 U4737 ( .A(n5051), .B(n5052), .Z(n5049));
  OR2 U4738 ( .A(n4319), .B(po013), .Z(n5052));
  OR2 U4739 ( .A(n5053), .B(po004), .Z(n5051));
  IV2 U4740 ( .A(po013), .Z(n5053));
  OR2 U4741 ( .A(n5054), .B(n5055), .Z(n5050));
  AN2 U4742 ( .A(po028), .B(n4013), .Z(n5055));
  AN2 U4743 ( .A(po040), .B(n5056), .Z(n5054));
  AN2 U4744 ( .A(n5057), .B(n5058), .Z(n5044));
  OR2 U4745 ( .A(n5059), .B(n5060), .Z(n5058));
  IV2 U4746 ( .A(n5061), .Z(n5059));
  OR2 U4747 ( .A(n5062), .B(n5061), .Z(n5057));
  OR2 U4748 ( .A(n5063), .B(n5064), .Z(n5061));
  AN2 U4749 ( .A(po064), .B(n4128), .Z(n5064));
  AN2 U4750 ( .A(po085), .B(n4133), .Z(n5063));
  IV2 U4751 ( .A(n5060), .Z(n5062));
  OR2 U4752 ( .A(n5065), .B(n5066), .Z(n5060));
  AN2 U4753 ( .A(po091), .B(n3265), .Z(n5066));
  AN2 U4754 ( .A(po103), .B(n4201), .Z(n5065));
  IV2 U4755 ( .A(n5067), .Z(po041));
  AN2 U4756 ( .A(n5068), .B(pi193), .Z(n5067));
  AN2 U4757 ( .A(pi057), .B(n5069), .Z(n5068));
  IV2 U4758 ( .A(pi037), .Z(n5069));
  OR2 U4759 ( .A(n5070), .B(n5071), .Z(po037));
  AN2 U4760 ( .A(n3021), .B(n5072), .Z(n5071));
  OR2 U4761 ( .A(n5073), .B(n5074), .Z(n5072));
  AN2 U4762 ( .A(n3018), .B(n5075), .Z(n5073));
  OR2 U4763 ( .A(n5076), .B(n5077), .Z(n5075));
  AN2 U4764 ( .A(n4663), .B(n3284), .Z(n5076));
  OR2 U4765 ( .A(n5078), .B(n5079), .Z(n4663));
  AN2 U4766 ( .A(n3064), .B(n3108), .Z(n5079));
  AN2 U4767 ( .A(n3173), .B(n3115), .Z(n5078));
  AN2 U4768 ( .A(n3083), .B(n5080), .Z(n5070));
  OR2 U4769 ( .A(n5081), .B(n5082), .Z(n5080));
  OR2 U4770 ( .A(n5083), .B(n5084), .Z(n5082));
  AN2 U4771 ( .A(po070), .B(n4327), .Z(n5084));
  OR2 U4772 ( .A(n5085), .B(n5086), .Z(n4327));
  OR2 U4773 ( .A(n5087), .B(n5088), .Z(n5086));
  AN2 U4774 ( .A(n3273), .B(n5089), .Z(n5088));
  IV2 U4775 ( .A(n3284), .Z(n3273));
  AN2 U4776 ( .A(n5090), .B(n3274), .Z(n5087));
  OR2 U4777 ( .A(n5091), .B(n3282), .Z(n5085));
  IV2 U4778 ( .A(n4666), .Z(n3282));
  AN2 U4779 ( .A(n5092), .B(n3199), .Z(n5083));
  OR2 U4780 ( .A(n5093), .B(n5094), .Z(n5092));
  OR2 U4781 ( .A(n5095), .B(n5096), .Z(n5094));
  AN2 U4782 ( .A(n5090), .B(po010), .Z(n5096));
  AN2 U4783 ( .A(n3037), .B(n3061), .Z(n5090));
  AN2 U4784 ( .A(n5097), .B(n5098), .Z(n5095));
  AN2 U4785 ( .A(n3037), .B(n5099), .Z(n5098));
  AN2 U4786 ( .A(n5100), .B(n3120), .Z(n5097));
  OR2 U4787 ( .A(n5101), .B(n3061), .Z(n3120));
  AN2 U4788 ( .A(n3106), .B(pi192), .Z(n3061));
  AN2 U4789 ( .A(po010), .B(pi192), .Z(n5101));
  AN2 U4790 ( .A(n3082), .B(pi192), .Z(n5093));
  IV2 U4791 ( .A(n3108), .Z(n3082));
  OR2 U4792 ( .A(pi033), .B(n3286), .Z(n3108));
  OR2 U4793 ( .A(n5102), .B(n5103), .Z(n5081));
  AN2 U4794 ( .A(n3015), .B(n5104), .Z(n5103));
  IV2 U4795 ( .A(n3018), .Z(n3015));
  AN2 U4796 ( .A(n5105), .B(n3205), .Z(n5102));
  OR2 U4797 ( .A(n5106), .B(n5107), .Z(n5105));
  OR2 U4798 ( .A(n5091), .B(n5108), .Z(n5107));
  AN2 U4799 ( .A(n5100), .B(n5109), .Z(n5108));
  OR2 U4800 ( .A(n5110), .B(n5111), .Z(n5109));
  AN2 U4801 ( .A(n5112), .B(n2925), .Z(n5111));
  AN2 U4802 ( .A(po010), .B(n5089), .Z(n5112));
  IV2 U4803 ( .A(n3100), .Z(n5089));
  AN2 U4804 ( .A(n5113), .B(n3080), .Z(n5110));
  AN2 U4805 ( .A(n2837), .B(po010), .Z(n3080));
  AN2 U4806 ( .A(n3112), .B(n5099), .Z(n5113));
  AN2 U4807 ( .A(n3065), .B(n5114), .Z(n5091));
  AN2 U4808 ( .A(n3112), .B(n3274), .Z(n5114));
  IV2 U4809 ( .A(n3280), .Z(n3274));
  AN2 U4810 ( .A(n2837), .B(n5115), .Z(n3065));
  AN2 U4811 ( .A(n3073), .B(n2837), .Z(n5106));
  IV2 U4812 ( .A(n3115), .Z(n3073));
  OR2 U4813 ( .A(pi141), .B(n3286), .Z(n3115));
  OR2 U4814 ( .A(n5116), .B(n5117), .Z(po034));
  OR2 U4815 ( .A(n5118), .B(n5119), .Z(n5117));
  AN2 U4816 ( .A(pi054), .B(n5120), .Z(n5119));
  AN2 U4817 ( .A(n5121), .B(n5122), .Z(n5118));
  AN2 U4818 ( .A(n5123), .B(n5124), .Z(n5122));
  OR2 U4819 ( .A(po085), .B(po064), .Z(n5124));
  OR2 U4820 ( .A(n4125), .B(n4133), .Z(n5123));
  AN2 U4821 ( .A(n4129), .B(n4128), .Z(n4125));
  AN2 U4822 ( .A(pi052), .B(n5125), .Z(n5121));
  AN2 U4823 ( .A(n5126), .B(n5127), .Z(n5116));
  OR2 U4824 ( .A(n4167), .B(n5128), .Z(n5127));
  OR2 U4825 ( .A(n5129), .B(n5130), .Z(n5128));
  AN2 U4826 ( .A(n5131), .B(po064), .Z(n5130));
  AN2 U4827 ( .A(pi054), .B(po085), .Z(n5131));
  AN2 U4828 ( .A(n4129), .B(n4133), .Z(n5129));
  OR2 U4829 ( .A(n5132), .B(n5133), .Z(po033));
  AN2 U4830 ( .A(n3371), .B(n5134), .Z(n5133));
  OR2 U4831 ( .A(n5135), .B(n5136), .Z(n5134));
  AN2 U4832 ( .A(n5137), .B(n3412), .Z(n5132));
  OR2 U4833 ( .A(n5138), .B(n5139), .Z(n5137));
  OR2 U4834 ( .A(n5140), .B(n5141), .Z(po030));
  AN2 U4835 ( .A(n5142), .B(pi192), .Z(n5141));
  OR2 U4836 ( .A(n5143), .B(n5144), .Z(n5142));
  AN2 U4837 ( .A(n2834), .B(n5145), .Z(n5144));
  OR2 U4838 ( .A(n5146), .B(n5147), .Z(n5145));
  AN2 U4839 ( .A(n2998), .B(n3847), .Z(n5147));
  AN2 U4840 ( .A(n5148), .B(n5149), .Z(n5146));
  OR2 U4841 ( .A(n2862), .B(n5150), .Z(n5149));
  OR2 U4842 ( .A(n2880), .B(n5151), .Z(n5150));
  AN2 U4843 ( .A(n2887), .B(n2901), .Z(n5151));
  AN2 U4844 ( .A(n2891), .B(n5152), .Z(n5148));
  IV2 U4845 ( .A(n5153), .Z(n5152));
  AN2 U4846 ( .A(n5154), .B(n2833), .Z(n5143));
  OR2 U4847 ( .A(n5155), .B(n5156), .Z(n5154));
  AN2 U4848 ( .A(n5157), .B(n5158), .Z(n5155));
  AN2 U4849 ( .A(n2930), .B(n2878), .Z(n5158));
  AN2 U4850 ( .A(n5159), .B(n2837), .Z(n5140));
  OR2 U4851 ( .A(n5160), .B(n5161), .Z(n5159));
  AN2 U4852 ( .A(n2846), .B(n5162), .Z(n5161));
  OR2 U4853 ( .A(n5163), .B(n5164), .Z(n5162));
  AN2 U4854 ( .A(n2998), .B(n5165), .Z(n5164));
  AN2 U4855 ( .A(n5166), .B(n5167), .Z(n5163));
  OR2 U4856 ( .A(n5168), .B(n5169), .Z(n5167));
  AN2 U4857 ( .A(n3222), .B(n2946), .Z(n5168));
  OR2 U4858 ( .A(n5170), .B(n2959), .Z(n3222));
  AN2 U4859 ( .A(n2982), .B(n2901), .Z(n2959));
  AN2 U4860 ( .A(po107), .B(n5171), .Z(n5170));
  IV2 U4861 ( .A(n2981), .Z(n5171));
  AN2 U4862 ( .A(pi081), .B(pi200), .Z(n2981));
  AN2 U4863 ( .A(n2947), .B(n5172), .Z(n5166));
  AN2 U4864 ( .A(n5173), .B(n2845), .Z(n5160));
  OR2 U4865 ( .A(n5174), .B(n5175), .Z(n5173));
  AN2 U4866 ( .A(n5157), .B(n5176), .Z(n5174));
  AN2 U4867 ( .A(n2908), .B(n2938), .Z(n5176));
  OR2 U4868 ( .A(pi081), .B(n2931), .Z(n2938));
  IV2 U4869 ( .A(n5169), .Z(n2908));
  AN2 U4870 ( .A(n2861), .B(pi200), .Z(n5157));
  OR2 U4871 ( .A(n5177), .B(n5178), .Z(po029));
  OR2 U4872 ( .A(n5179), .B(n5180), .Z(n5178));
  AN2 U4873 ( .A(n5181), .B(n4313), .Z(n5180));
  AN2 U4874 ( .A(n3945), .B(n5182), .Z(n5179));
  OR2 U4875 ( .A(n5183), .B(n5184), .Z(n5182));
  OR2 U4876 ( .A(n5185), .B(n5186), .Z(n5184));
  AN2 U4877 ( .A(n5187), .B(pi186), .Z(n5186));
  OR2 U4878 ( .A(n5188), .B(n5189), .Z(n5187));
  AN2 U4879 ( .A(n5190), .B(n5191), .Z(n5189));
  AN2 U4880 ( .A(n5192), .B(pi124), .Z(n5188));
  IV2 U4881 ( .A(n5190), .Z(n5192));
  AN2 U4882 ( .A(n5193), .B(n5194), .Z(n5185));
  OR2 U4883 ( .A(n5195), .B(n5196), .Z(n5193));
  AN2 U4884 ( .A(n5190), .B(pi124), .Z(n5196));
  OR2 U4885 ( .A(n5197), .B(n5198), .Z(n5190));
  AN2 U4886 ( .A(n5199), .B(n5200), .Z(n5198));
  AN2 U4887 ( .A(n5201), .B(pi109), .Z(n5197));
  IV2 U4888 ( .A(n5199), .Z(n5201));
  AN2 U4889 ( .A(n5202), .B(n5191), .Z(n5195));
  OR2 U4890 ( .A(n5203), .B(n5204), .Z(n5202));
  AN2 U4891 ( .A(n5199), .B(pi109), .Z(n5204));
  OR2 U4892 ( .A(n5205), .B(n5206), .Z(n5199));
  AN2 U4893 ( .A(n5207), .B(n5208), .Z(n5206));
  AN2 U4894 ( .A(n5181), .B(pi055), .Z(n5205));
  AN2 U4895 ( .A(n5209), .B(n5200), .Z(n5203));
  AN2 U4896 ( .A(pi055), .B(n5207), .Z(n5209));
  AN2 U4897 ( .A(n5210), .B(n5211), .Z(n5183));
  OR2 U4898 ( .A(n5212), .B(n5213), .Z(n5211));
  IV2 U4899 ( .A(n5214), .Z(n5210));
  AN2 U4900 ( .A(n5213), .B(n5212), .Z(n5214));
  OR2 U4901 ( .A(n5215), .B(n5216), .Z(n5212));
  IV2 U4902 ( .A(n5217), .Z(n5216));
  OR2 U4903 ( .A(n5218), .B(pi006), .Z(n5217));
  AN2 U4904 ( .A(n5218), .B(pi006), .Z(n5215));
  AN2 U4905 ( .A(n5219), .B(n5220), .Z(n5218));
  OR2 U4906 ( .A(n5221), .B(pi061), .Z(n5220));
  IV2 U4907 ( .A(pi051), .Z(n5221));
  OR2 U4908 ( .A(n5222), .B(pi051), .Z(n5219));
  IV2 U4909 ( .A(pi061), .Z(n5222));
  AN2 U4910 ( .A(n5223), .B(n5224), .Z(n5213));
  IV2 U4911 ( .A(n5225), .Z(n5224));
  AN2 U4912 ( .A(n5226), .B(n5227), .Z(n5225));
  OR2 U4913 ( .A(n5227), .B(n5226), .Z(n5223));
  OR2 U4914 ( .A(n5228), .B(n5229), .Z(n5226));
  AN2 U4915 ( .A(pi093), .B(n5230), .Z(n5229));
  IV2 U4916 ( .A(n5231), .Z(n5228));
  OR2 U4917 ( .A(n5230), .B(pi093), .Z(n5231));
  IV2 U4918 ( .A(pi122), .Z(n5230));
  AN2 U4919 ( .A(n5232), .B(n5233), .Z(n5227));
  IV2 U4920 ( .A(n5234), .Z(n5233));
  AN2 U4921 ( .A(pi134), .B(n5235), .Z(n5234));
  OR2 U4922 ( .A(n5235), .B(pi134), .Z(n5232));
  IV2 U4923 ( .A(pi198), .Z(n5235));
  OR2 U4924 ( .A(n5236), .B(n5237), .Z(n5177));
  AN2 U4925 ( .A(n5238), .B(n2837), .Z(n5237));
  OR2 U4926 ( .A(n5239), .B(n5240), .Z(n5238));
  AN2 U4927 ( .A(n5241), .B(n5242), .Z(n5240));
  OR2 U4928 ( .A(n3809), .B(n5243), .Z(n5242));
  IV2 U4929 ( .A(n3812), .Z(n3809));
  OR2 U4930 ( .A(n5244), .B(n3812), .Z(n5241));
  AN2 U4931 ( .A(n5245), .B(n5246), .Z(n3812));
  IV2 U4932 ( .A(n5247), .Z(n5246));
  AN2 U4933 ( .A(n5248), .B(n5249), .Z(n5247));
  OR2 U4934 ( .A(n5249), .B(n5248), .Z(n5245));
  OR2 U4935 ( .A(n5250), .B(n5251), .Z(n5248));
  AN2 U4936 ( .A(pi040), .B(n5252), .Z(n5251));
  IV2 U4937 ( .A(pi095), .Z(n5252));
  AN2 U4938 ( .A(pi095), .B(n4735), .Z(n5250));
  AN2 U4939 ( .A(n5253), .B(n5254), .Z(n5249));
  OR2 U4940 ( .A(n4747), .B(pi156), .Z(n5254));
  IV2 U4941 ( .A(pi151), .Z(n4747));
  OR2 U4942 ( .A(n4648), .B(pi151), .Z(n5253));
  AN2 U4943 ( .A(n5255), .B(n5256), .Z(n5239));
  OR2 U4944 ( .A(n3815), .B(n5257), .Z(n5256));
  OR2 U4945 ( .A(n5258), .B(n3818), .Z(n5255));
  IV2 U4946 ( .A(n3815), .Z(n3818));
  OR2 U4947 ( .A(n5259), .B(n5260), .Z(n3815));
  AN2 U4948 ( .A(n5261), .B(n5262), .Z(n5260));
  IV2 U4949 ( .A(n5263), .Z(n5259));
  OR2 U4950 ( .A(n5262), .B(n5261), .Z(n5263));
  OR2 U4951 ( .A(n5264), .B(n5265), .Z(n5261));
  AN2 U4952 ( .A(pi128), .B(n3177), .Z(n5265));
  AN2 U4953 ( .A(pi141), .B(n3205), .Z(n5264));
  AN2 U4954 ( .A(n5266), .B(n5267), .Z(n5262));
  OR2 U4955 ( .A(n5115), .B(pi185), .Z(n5267));
  OR2 U4956 ( .A(n5268), .B(pi174), .Z(n5266));
  IV2 U4957 ( .A(pi185), .Z(n5268));
  AN2 U4958 ( .A(pi192), .B(n5269), .Z(n5236));
  OR2 U4959 ( .A(n5270), .B(n5271), .Z(n5269));
  OR2 U4960 ( .A(n5272), .B(n5273), .Z(n5271));
  AN2 U4961 ( .A(n5274), .B(n5275), .Z(n5273));
  IV2 U4962 ( .A(n5276), .Z(n5275));
  AN2 U4963 ( .A(n5277), .B(n5278), .Z(n5276));
  OR2 U4964 ( .A(n5278), .B(n5277), .Z(n5274));
  AN2 U4965 ( .A(n5279), .B(n5280), .Z(n5277));
  OR2 U4966 ( .A(n5243), .B(pi036), .Z(n5280));
  IV2 U4967 ( .A(n5244), .Z(n5243));
  OR2 U4968 ( .A(n5244), .B(n5281), .Z(n5279));
  IV2 U4969 ( .A(pi036), .Z(n5281));
  OR2 U4970 ( .A(n3871), .B(n5282), .Z(n5244));
  AN2 U4971 ( .A(n5283), .B(pi192), .Z(n5282));
  OR2 U4972 ( .A(n5284), .B(n5285), .Z(n5283));
  AN2 U4973 ( .A(n5286), .B(n5287), .Z(n5285));
  IV2 U4974 ( .A(n5288), .Z(n5284));
  OR2 U4975 ( .A(n5287), .B(n5286), .Z(n5288));
  OR2 U4976 ( .A(n5289), .B(n5290), .Z(n5286));
  IV2 U4977 ( .A(n5291), .Z(n5290));
  OR2 U4978 ( .A(n5292), .B(pi017), .Z(n5291));
  AN2 U4979 ( .A(pi017), .B(n5292), .Z(n5289));
  AN2 U4980 ( .A(n5293), .B(n5294), .Z(n5292));
  OR2 U4981 ( .A(n5295), .B(pi083), .Z(n5294));
  IV2 U4982 ( .A(pi027), .Z(n5295));
  OR2 U4983 ( .A(n5296), .B(pi027), .Z(n5293));
  IV2 U4984 ( .A(pi083), .Z(n5296));
  AN2 U4985 ( .A(n5297), .B(n5298), .Z(n5287));
  OR2 U4986 ( .A(n5299), .B(pi089), .Z(n5298));
  IV2 U4987 ( .A(n5300), .Z(n5297));
  AN2 U4988 ( .A(n5299), .B(pi089), .Z(n5300));
  AN2 U4989 ( .A(n5301), .B(n5302), .Z(n5299));
  OR2 U4990 ( .A(n5303), .B(pi162), .Z(n5302));
  OR2 U4991 ( .A(n5304), .B(pi140), .Z(n5301));
  IV2 U4992 ( .A(pi162), .Z(n5304));
  AN2 U4993 ( .A(n5305), .B(n2837), .Z(n3871));
  OR2 U4994 ( .A(n5306), .B(n5307), .Z(n5305));
  AN2 U4995 ( .A(n5308), .B(n5309), .Z(n5307));
  IV2 U4996 ( .A(n5310), .Z(n5306));
  OR2 U4997 ( .A(n5309), .B(n5308), .Z(n5310));
  OR2 U4998 ( .A(n5311), .B(n5312), .Z(n5308));
  IV2 U4999 ( .A(n5313), .Z(n5312));
  OR2 U5000 ( .A(n5314), .B(pi064), .Z(n5313));
  AN2 U5001 ( .A(pi064), .B(n5314), .Z(n5311));
  AN2 U5002 ( .A(n5315), .B(n5316), .Z(n5314));
  OR2 U5003 ( .A(n4077), .B(pi108), .Z(n5316));
  OR2 U5004 ( .A(n5317), .B(pi076), .Z(n5315));
  IV2 U5005 ( .A(pi108), .Z(n5317));
  AN2 U5006 ( .A(n5318), .B(n5319), .Z(n5309));
  OR2 U5007 ( .A(n5320), .B(pi114), .Z(n5319));
  IV2 U5008 ( .A(n5321), .Z(n5320));
  OR2 U5009 ( .A(n5321), .B(n5322), .Z(n5318));
  OR2 U5010 ( .A(n5323), .B(n5324), .Z(n5321));
  AN2 U5011 ( .A(pi160), .B(n4074), .Z(n5324));
  AN2 U5012 ( .A(pi170), .B(n4358), .Z(n5323));
  OR2 U5013 ( .A(n5325), .B(n5326), .Z(n5278));
  IV2 U5014 ( .A(n5327), .Z(n5326));
  OR2 U5015 ( .A(n5328), .B(pi101), .Z(n5327));
  AN2 U5016 ( .A(n5328), .B(pi101), .Z(n5325));
  AN2 U5017 ( .A(n5329), .B(n5330), .Z(n5328));
  OR2 U5018 ( .A(n5331), .B(pi205), .Z(n5330));
  OR2 U5019 ( .A(n5332), .B(pi168), .Z(n5329));
  IV2 U5020 ( .A(pi205), .Z(n5332));
  AN2 U5021 ( .A(n5333), .B(n5334), .Z(n5272));
  AN2 U5022 ( .A(n5335), .B(n5200), .Z(n5334));
  IV2 U5023 ( .A(pi109), .Z(n5200));
  AN2 U5024 ( .A(n5191), .B(n5194), .Z(n5335));
  IV2 U5025 ( .A(pi186), .Z(n5194));
  IV2 U5026 ( .A(pi124), .Z(n5191));
  AN2 U5027 ( .A(n5181), .B(n5208), .Z(n5333));
  IV2 U5028 ( .A(pi055), .Z(n5208));
  IV2 U5029 ( .A(n5207), .Z(n5181));
  OR2 U5030 ( .A(n3977), .B(n5336), .Z(n5207));
  AN2 U5031 ( .A(n5337), .B(pi192), .Z(n5336));
  OR2 U5032 ( .A(n5338), .B(n5339), .Z(n5337));
  AN2 U5033 ( .A(n5340), .B(n5341), .Z(n5339));
  IV2 U5034 ( .A(n5342), .Z(n5338));
  OR2 U5035 ( .A(n5341), .B(n5340), .Z(n5342));
  OR2 U5036 ( .A(n5343), .B(n5344), .Z(n5340));
  IV2 U5037 ( .A(n5345), .Z(n5344));
  OR2 U5038 ( .A(n5346), .B(n5347), .Z(n5345));
  AN2 U5039 ( .A(n5346), .B(n5347), .Z(n5343));
  AN2 U5040 ( .A(n5348), .B(n5349), .Z(n5346));
  OR2 U5041 ( .A(n5350), .B(pi099), .Z(n5349));
  OR2 U5042 ( .A(n5351), .B(pi018), .Z(n5348));
  IV2 U5043 ( .A(pi099), .Z(n5351));
  AN2 U5044 ( .A(n5352), .B(n5353), .Z(n5341));
  OR2 U5045 ( .A(n5354), .B(pi150), .Z(n5353));
  IV2 U5046 ( .A(n5355), .Z(n5352));
  AN2 U5047 ( .A(pi150), .B(n5354), .Z(n5355));
  AN2 U5048 ( .A(n5356), .B(n5357), .Z(n5354));
  OR2 U5049 ( .A(n5358), .B(pi180), .Z(n5357));
  OR2 U5050 ( .A(n5359), .B(pi172), .Z(n5356));
  IV2 U5051 ( .A(pi180), .Z(n5359));
  AN2 U5052 ( .A(n5360), .B(n2837), .Z(n3977));
  AN2 U5053 ( .A(n5361), .B(n5362), .Z(n5360));
  IV2 U5054 ( .A(n5363), .Z(n5362));
  AN2 U5055 ( .A(n5364), .B(n5365), .Z(n5363));
  OR2 U5056 ( .A(n5365), .B(n5364), .Z(n5361));
  OR2 U5057 ( .A(n5366), .B(n5367), .Z(n5364));
  AN2 U5058 ( .A(n5368), .B(n3261), .Z(n5367));
  AN2 U5059 ( .A(n5369), .B(n3321), .Z(n5366));
  IV2 U5060 ( .A(n5368), .Z(n5369));
  OR2 U5061 ( .A(n5370), .B(n5371), .Z(n5368));
  AN2 U5062 ( .A(pi003), .B(n5372), .Z(n5371));
  AN2 U5063 ( .A(pi130), .B(n3597), .Z(n5370));
  AN2 U5064 ( .A(n5373), .B(n5374), .Z(n5365));
  OR2 U5065 ( .A(n5375), .B(pi142), .Z(n5374));
  IV2 U5066 ( .A(n5376), .Z(n5375));
  OR2 U5067 ( .A(n5376), .B(n4440), .Z(n5373));
  OR2 U5068 ( .A(n5377), .B(n5378), .Z(n5376));
  AN2 U5069 ( .A(pi177), .B(n5379), .Z(n5378));
  AN2 U5070 ( .A(pi195), .B(n5380), .Z(n5377));
  IV2 U5071 ( .A(pi177), .Z(n5380));
  AN2 U5072 ( .A(n5381), .B(n5382), .Z(n5270));
  IV2 U5073 ( .A(n5383), .Z(n5382));
  AN2 U5074 ( .A(n5384), .B(n5385), .Z(n5383));
  OR2 U5075 ( .A(n5385), .B(n5384), .Z(n5381));
  AN2 U5076 ( .A(n5386), .B(n5387), .Z(n5384));
  OR2 U5077 ( .A(n5257), .B(pi001), .Z(n5387));
  IV2 U5078 ( .A(n5258), .Z(n5257));
  OR2 U5079 ( .A(n5258), .B(n5388), .Z(n5386));
  IV2 U5080 ( .A(pi001), .Z(n5388));
  OR2 U5081 ( .A(n3831), .B(n5389), .Z(n5258));
  AN2 U5082 ( .A(n5390), .B(pi192), .Z(n5389));
  OR2 U5083 ( .A(n5391), .B(n5392), .Z(n5390));
  AN2 U5084 ( .A(n5393), .B(n5394), .Z(n5392));
  IV2 U5085 ( .A(n5395), .Z(n5391));
  OR2 U5086 ( .A(n5394), .B(n5393), .Z(n5395));
  OR2 U5087 ( .A(n5396), .B(n5397), .Z(n5393));
  IV2 U5088 ( .A(n5398), .Z(n5397));
  OR2 U5089 ( .A(n5399), .B(pi038), .Z(n5398));
  AN2 U5090 ( .A(pi038), .B(n5399), .Z(n5396));
  AN2 U5091 ( .A(n5400), .B(n5401), .Z(n5399));
  OR2 U5092 ( .A(n5402), .B(pi103), .Z(n5401));
  IV2 U5093 ( .A(pi053), .Z(n5402));
  OR2 U5094 ( .A(n5403), .B(pi053), .Z(n5400));
  IV2 U5095 ( .A(pi103), .Z(n5403));
  AN2 U5096 ( .A(n5404), .B(n5405), .Z(n5394));
  OR2 U5097 ( .A(n5406), .B(pi121), .Z(n5405));
  IV2 U5098 ( .A(n5407), .Z(n5404));
  AN2 U5099 ( .A(n5406), .B(pi121), .Z(n5407));
  AN2 U5100 ( .A(n5408), .B(n5409), .Z(n5406));
  OR2 U5101 ( .A(n5410), .B(pi184), .Z(n5409));
  IV2 U5102 ( .A(pi149), .Z(n5410));
  OR2 U5103 ( .A(n5411), .B(pi149), .Z(n5408));
  IV2 U5104 ( .A(pi184), .Z(n5411));
  AN2 U5105 ( .A(n5412), .B(n2837), .Z(n3831));
  OR2 U5106 ( .A(n5413), .B(n5414), .Z(n5412));
  IV2 U5107 ( .A(n5415), .Z(n5414));
  OR2 U5108 ( .A(n5416), .B(n5417), .Z(n5415));
  AN2 U5109 ( .A(n5417), .B(n5416), .Z(n5413));
  AN2 U5110 ( .A(n5418), .B(n5419), .Z(n5416));
  OR2 U5111 ( .A(n5420), .B(pi081), .Z(n5419));
  IV2 U5112 ( .A(n5421), .Z(n5420));
  OR2 U5113 ( .A(n5421), .B(n2982), .Z(n5418));
  OR2 U5114 ( .A(n5422), .B(n5423), .Z(n5421));
  AN2 U5115 ( .A(pi082), .B(n5424), .Z(n5423));
  IV2 U5116 ( .A(pi092), .Z(n5424));
  AN2 U5117 ( .A(pi092), .B(n2957), .Z(n5422));
  OR2 U5118 ( .A(n5425), .B(n5426), .Z(n5417));
  AN2 U5119 ( .A(n5427), .B(n5165), .Z(n5426));
  AN2 U5120 ( .A(n5428), .B(pi107), .Z(n5425));
  IV2 U5121 ( .A(n5427), .Z(n5428));
  OR2 U5122 ( .A(n5429), .B(n5430), .Z(n5427));
  AN2 U5123 ( .A(pi201), .B(n5431), .Z(n5430));
  AN2 U5124 ( .A(pi206), .B(n3141), .Z(n5429));
  OR2 U5125 ( .A(n5432), .B(n5433), .Z(n5385));
  IV2 U5126 ( .A(n5434), .Z(n5433));
  OR2 U5127 ( .A(n5435), .B(pi059), .Z(n5434));
  AN2 U5128 ( .A(n5435), .B(pi059), .Z(n5432));
  AN2 U5129 ( .A(n5436), .B(n5437), .Z(n5435));
  OR2 U5130 ( .A(n5438), .B(pi197), .Z(n5437));
  IV2 U5131 ( .A(pi131), .Z(n5438));
  OR2 U5132 ( .A(n5439), .B(pi131), .Z(n5436));
  OR2 U5133 ( .A(n5440), .B(n5441), .Z(po026));
  AN2 U5134 ( .A(n3355), .B(n5442), .Z(n5441));
  OR2 U5135 ( .A(n5443), .B(n5444), .Z(n5442));
  OR2 U5136 ( .A(n5445), .B(n5446), .Z(n5444));
  AN2 U5137 ( .A(po036), .B(n5447), .Z(n5446));
  OR2 U5138 ( .A(n4418), .B(n5448), .Z(n5447));
  AN2 U5139 ( .A(n5449), .B(n3236), .Z(n5445));
  AN2 U5140 ( .A(n5450), .B(n5451), .Z(n5449));
  OR2 U5141 ( .A(n5452), .B(n2837), .Z(n5451));
  OR2 U5142 ( .A(pi192), .B(n5453), .Z(n5450));
  AN2 U5143 ( .A(n4418), .B(n5448), .Z(n5443));
  AN2 U5144 ( .A(n3352), .B(n5454), .Z(n5440));
  IV2 U5145 ( .A(n5455), .Z(po022));
  AN2 U5146 ( .A(n5456), .B(n5457), .Z(n5455));
  AN2 U5147 ( .A(pi074), .B(pi046), .Z(n5457));
  AN2 U5148 ( .A(pi178), .B(pi113), .Z(n5456));
  OR2 U5149 ( .A(n5458), .B(n5459), .Z(po019));
  AN2 U5150 ( .A(n4478), .B(n5460), .Z(n5459));
  OR2 U5151 ( .A(n5461), .B(n4511), .Z(n5460));
  OR2 U5152 ( .A(n5462), .B(n5463), .Z(n4511));
  OR2 U5153 ( .A(n5464), .B(n5465), .Z(n5463));
  AN2 U5154 ( .A(n5466), .B(pi192), .Z(n5465));
  AN2 U5155 ( .A(n5467), .B(n2837), .Z(n5464));
  AN2 U5156 ( .A(n4475), .B(n5468), .Z(n5458));
  OR2 U5157 ( .A(n5469), .B(n5470), .Z(n5468));
  OR2 U5158 ( .A(n5471), .B(n4509), .Z(n5470));
  OR2 U5159 ( .A(n5472), .B(n5473), .Z(n4509));
  OR2 U5160 ( .A(n5474), .B(n5475), .Z(n5473));
  AN2 U5161 ( .A(n5476), .B(n4078), .Z(n5475));
  AN2 U5162 ( .A(n5477), .B(n5322), .Z(n5476));
  AN2 U5163 ( .A(n5478), .B(n4551), .Z(n5472));
  IV2 U5164 ( .A(n4544), .Z(n4551));
  OR2 U5165 ( .A(n4561), .B(n4066), .Z(n4544));
  AN2 U5166 ( .A(pi192), .B(n3901), .Z(n5478));
  AN2 U5167 ( .A(po102), .B(n4347), .Z(n5471));
  OR2 U5168 ( .A(n5479), .B(n4524), .Z(n4347));
  AN2 U5169 ( .A(n5480), .B(n4078), .Z(n4524));
  IV2 U5170 ( .A(n4066), .Z(n4078));
  AN2 U5171 ( .A(n4521), .B(n4072), .Z(n5479));
  OR2 U5172 ( .A(n5481), .B(n5482), .Z(n4521));
  AN2 U5173 ( .A(po059), .B(n5480), .Z(n5482));
  OR2 U5174 ( .A(n5483), .B(po024), .Z(n5480));
  AN2 U5175 ( .A(n5477), .B(n4074), .Z(n5481));
  OR2 U5176 ( .A(n5484), .B(n5485), .Z(n5469));
  AN2 U5177 ( .A(n4517), .B(n3780), .Z(n5485));
  OR2 U5178 ( .A(n5486), .B(n5487), .Z(n4517));
  AN2 U5179 ( .A(n4356), .B(n5488), .Z(n5487));
  AN2 U5180 ( .A(n4076), .B(n5489), .Z(n4356));
  AN2 U5181 ( .A(n4077), .B(n4578), .Z(n5489));
  AN2 U5182 ( .A(n5490), .B(n4543), .Z(n5486));
  AN2 U5183 ( .A(n4348), .B(n4353), .Z(n4543));
  AN2 U5184 ( .A(n3890), .B(n5491), .Z(n5490));
  AN2 U5185 ( .A(n4512), .B(n4072), .Z(n5484));
  OR2 U5186 ( .A(n5492), .B(n3773), .Z(n4072));
  AN2 U5187 ( .A(po025), .B(n3780), .Z(n5492));
  IV2 U5188 ( .A(n4087), .Z(n3780));
  OR2 U5189 ( .A(n5493), .B(n5494), .Z(n4512));
  OR2 U5190 ( .A(n5495), .B(n5496), .Z(n5494));
  AN2 U5191 ( .A(n5497), .B(pi192), .Z(n5496));
  AN2 U5192 ( .A(n5498), .B(n4348), .Z(n5497));
  OR2 U5193 ( .A(n5499), .B(n5500), .Z(n5498));
  AN2 U5194 ( .A(po102), .B(n3880), .Z(n5500));
  AN2 U5195 ( .A(n4353), .B(n3901), .Z(n5499));
  AN2 U5196 ( .A(n5501), .B(n4076), .Z(n5495));
  AN2 U5197 ( .A(n5488), .B(n4358), .Z(n5501));
  AN2 U5198 ( .A(n5502), .B(n4076), .Z(n5493));
  AN2 U5199 ( .A(n2837), .B(n5503), .Z(n4076));
  AN2 U5200 ( .A(po024), .B(n5322), .Z(n5502));
  OR2 U5201 ( .A(n5504), .B(n5505), .Z(po074));
  AN2 U5202 ( .A(n5506), .B(n5507), .Z(n5505));
  OR2 U5203 ( .A(n4167), .B(n5508), .Z(n5507));
  OR2 U5204 ( .A(pi054), .B(n5509), .Z(n5508));
  AN2 U5205 ( .A(pi025), .B(pi146), .Z(n5509));
  OR2 U5206 ( .A(n5510), .B(n5511), .Z(n5506));
  OR2 U5207 ( .A(n5512), .B(n5513), .Z(n5511));
  AN2 U5208 ( .A(n3926), .B(n5514), .Z(n5513));
  OR2 U5209 ( .A(n5515), .B(n5516), .Z(n5514));
  OR2 U5210 ( .A(n5517), .B(n5518), .Z(n5516));
  OR2 U5211 ( .A(pi056), .B(pi035), .Z(n5518));
  OR2 U5212 ( .A(pi100), .B(n5519), .Z(n5515));
  OR2 U5213 ( .A(pi190), .B(pi126), .Z(n5519));
  AN2 U5214 ( .A(n5520), .B(n4319), .Z(n5512));
  OR2 U5215 ( .A(n5521), .B(n5522), .Z(n5520));
  AN2 U5216 ( .A(pi198), .B(n3945), .Z(n5522));
  AN2 U5217 ( .A(n5523), .B(n5524), .Z(n5521));
  AN2 U5218 ( .A(n5525), .B(n5517), .Z(n5524));
  AN2 U5219 ( .A(n5056), .B(n4201), .Z(n5525));
  AN2 U5220 ( .A(n4391), .B(pi192), .Z(n5523));
  OR2 U5221 ( .A(n5526), .B(n5527), .Z(n5510));
  AN2 U5222 ( .A(n5528), .B(n5529), .Z(n5527));
  OR2 U5223 ( .A(pi198), .B(n4319), .Z(n5529));
  OR2 U5224 ( .A(n5530), .B(n5531), .Z(n5528));
  AN2 U5225 ( .A(n3945), .B(n5532), .Z(n5531));
  OR2 U5226 ( .A(n5533), .B(n5534), .Z(n5532));
  AN2 U5227 ( .A(pi061), .B(n4013), .Z(n5534));
  AN2 U5228 ( .A(n5535), .B(pi134), .Z(n5533));
  AN2 U5229 ( .A(n5536), .B(n4201), .Z(n5535));
  AN2 U5230 ( .A(n5537), .B(n5538), .Z(n5530));
  AN2 U5231 ( .A(n5536), .B(n3261), .Z(n5538));
  OR2 U5232 ( .A(pi061), .B(n4013), .Z(n5536));
  AN2 U5233 ( .A(n5539), .B(n5540), .Z(n5537));
  OR2 U5234 ( .A(pi134), .B(n4201), .Z(n5540));
  OR2 U5235 ( .A(n5541), .B(n5542), .Z(n5539));
  AN2 U5236 ( .A(n5543), .B(n5517), .Z(n5542));
  AN2 U5237 ( .A(pi192), .B(n5544), .Z(n5541));
  OR2 U5238 ( .A(n5545), .B(n5546), .Z(n5544));
  AN2 U5239 ( .A(pi006), .B(n3265), .Z(n5546));
  AN2 U5240 ( .A(n5543), .B(n5056), .Z(n5545));
  OR2 U5241 ( .A(pi006), .B(n3265), .Z(n5543));
  AN2 U5242 ( .A(n5547), .B(n5548), .Z(n5526));
  AN2 U5243 ( .A(n5549), .B(n5550), .Z(n5548));
  AN2 U5244 ( .A(n5517), .B(n2837), .Z(n5550));
  OR2 U5245 ( .A(n5551), .B(n5552), .Z(n5517));
  OR2 U5246 ( .A(n5553), .B(n5554), .Z(n5552));
  AN2 U5247 ( .A(n3945), .B(n5555), .Z(n5554));
  OR2 U5248 ( .A(n5556), .B(n5557), .Z(n5555));
  OR2 U5249 ( .A(n5558), .B(n5559), .Z(n5557));
  AN2 U5250 ( .A(n5560), .B(n3380), .Z(n5559));
  AN2 U5251 ( .A(n5561), .B(n5562), .Z(n5558));
  OR2 U5252 ( .A(n5563), .B(n5564), .Z(n5561));
  AN2 U5253 ( .A(pi055), .B(n3512), .Z(n5564));
  AN2 U5254 ( .A(n5565), .B(pi124), .Z(n5563));
  AN2 U5255 ( .A(n5566), .B(n3363), .Z(n5565));
  AN2 U5256 ( .A(pi109), .B(n4975), .Z(n5556));
  AN2 U5257 ( .A(n5567), .B(n5568), .Z(n5553));
  OR2 U5258 ( .A(n5569), .B(n5570), .Z(n5568));
  OR2 U5259 ( .A(n5571), .B(n5572), .Z(n5570));
  AN2 U5260 ( .A(n5573), .B(n5566), .Z(n5572));
  OR2 U5261 ( .A(pi055), .B(n3512), .Z(n5566));
  AN2 U5262 ( .A(n5574), .B(n3261), .Z(n5573));
  OR2 U5263 ( .A(n5575), .B(n5576), .Z(n5574));
  AN2 U5264 ( .A(pi124), .B(n5562), .Z(n5576));
  OR2 U5265 ( .A(n5577), .B(n5560), .Z(n5562));
  AN2 U5266 ( .A(n5578), .B(n3380), .Z(n5577));
  AN2 U5267 ( .A(n5579), .B(n3363), .Z(n5575));
  OR2 U5268 ( .A(n5580), .B(n5560), .Z(n5579));
  AN2 U5269 ( .A(n5578), .B(pi186), .Z(n5560));
  OR2 U5270 ( .A(pi109), .B(n4975), .Z(n5578));
  AN2 U5271 ( .A(pi109), .B(n3380), .Z(n5580));
  AN2 U5272 ( .A(n5581), .B(n5582), .Z(n5571));
  AN2 U5273 ( .A(n4975), .B(n3380), .Z(n5582));
  AN2 U5274 ( .A(n5583), .B(n3363), .Z(n5581));
  OR2 U5275 ( .A(n5584), .B(n5585), .Z(n5583));
  AN2 U5276 ( .A(pi192), .B(n3512), .Z(n5585));
  AN2 U5277 ( .A(pi055), .B(n3261), .Z(n5584));
  OR2 U5278 ( .A(n3926), .B(n5586), .Z(n5569));
  AN2 U5279 ( .A(n5587), .B(n5588), .Z(n5586));
  AN2 U5280 ( .A(n5589), .B(pi110), .Z(n5588));
  AN2 U5281 ( .A(pi167), .B(n2837), .Z(n5589));
  AN2 U5282 ( .A(pi019), .B(pi085), .Z(n5587));
  AN2 U5283 ( .A(n5590), .B(n5591), .Z(n5567));
  OR2 U5284 ( .A(pi192), .B(n5592), .Z(n5591));
  AN2 U5285 ( .A(n5593), .B(n5594), .Z(n5592));
  OR2 U5286 ( .A(pi164), .B(n3261), .Z(n5594));
  OR2 U5287 ( .A(n5595), .B(n5596), .Z(n5593));
  OR2 U5288 ( .A(n5597), .B(n5598), .Z(n5596));
  AN2 U5289 ( .A(n5599), .B(pi024), .Z(n5598));
  AN2 U5290 ( .A(pi195), .B(n5600), .Z(n5597));
  OR2 U5291 ( .A(n5601), .B(n5599), .Z(n5600));
  AN2 U5292 ( .A(n5602), .B(n5603), .Z(n5599));
  IV2 U5293 ( .A(n5604), .Z(n5603));
  AN2 U5294 ( .A(n5605), .B(n5606), .Z(n5604));
  OR2 U5295 ( .A(n5607), .B(n5608), .Z(n5606));
  AN2 U5296 ( .A(n5609), .B(n5610), .Z(n5608));
  OR2 U5297 ( .A(n5611), .B(n4961), .Z(n5610));
  IV2 U5298 ( .A(pi030), .Z(n4961));
  AN2 U5299 ( .A(n5612), .B(n3597), .Z(n5611));
  OR2 U5300 ( .A(n5612), .B(n3597), .Z(n5609));
  AN2 U5301 ( .A(n4969), .B(n4440), .Z(n5607));
  OR2 U5302 ( .A(n4440), .B(n4969), .Z(n5605));
  IV2 U5303 ( .A(pi159), .Z(n4969));
  AN2 U5304 ( .A(pi024), .B(n5602), .Z(n5601));
  OR2 U5305 ( .A(pi087), .B(pi130), .Z(n5602));
  AN2 U5306 ( .A(pi087), .B(pi130), .Z(n5595));
  OR2 U5307 ( .A(n2837), .B(n5613), .Z(n5590));
  OR2 U5308 ( .A(n5614), .B(n5615), .Z(n5613));
  AN2 U5309 ( .A(n5347), .B(n5616), .Z(n5615));
  AN2 U5310 ( .A(n5617), .B(n4943), .Z(n5614));
  OR2 U5311 ( .A(n5347), .B(n5616), .Z(n5617));
  OR2 U5312 ( .A(n5618), .B(n5619), .Z(n5616));
  OR2 U5313 ( .A(n5620), .B(n5621), .Z(n5619));
  AN2 U5314 ( .A(n5622), .B(pi099), .Z(n5621));
  AN2 U5315 ( .A(n5623), .B(n4937), .Z(n5620));
  OR2 U5316 ( .A(n5624), .B(n5622), .Z(n5623));
  AN2 U5317 ( .A(n5625), .B(n5626), .Z(n5622));
  IV2 U5318 ( .A(n5627), .Z(n5626));
  AN2 U5319 ( .A(n5628), .B(n5629), .Z(n5627));
  OR2 U5320 ( .A(n5630), .B(n5631), .Z(n5629));
  AN2 U5321 ( .A(n5632), .B(n5633), .Z(n5631));
  OR2 U5322 ( .A(po011), .B(n5634), .Z(n5633));
  AN2 U5323 ( .A(n5612), .B(n5358), .Z(n5634));
  OR2 U5324 ( .A(n5612), .B(n5358), .Z(n5632));
  IV2 U5325 ( .A(pi172), .Z(n5358));
  IV2 U5326 ( .A(po062), .Z(n5612));
  OR2 U5327 ( .A(n5635), .B(n5636), .Z(po062));
  AN2 U5328 ( .A(n5637), .B(n2837), .Z(n5636));
  OR2 U5329 ( .A(n5638), .B(n5639), .Z(n5637));
  AN2 U5330 ( .A(pi020), .B(pi095), .Z(n5639));
  AN2 U5331 ( .A(n5640), .B(n5641), .Z(n5638));
  OR2 U5332 ( .A(pi020), .B(pi095), .Z(n5641));
  OR2 U5333 ( .A(n5642), .B(n5643), .Z(n5640));
  AN2 U5334 ( .A(pi151), .B(n5644), .Z(n5643));
  AN2 U5335 ( .A(pi153), .B(n5645), .Z(n5642));
  OR2 U5336 ( .A(pi151), .B(n5644), .Z(n5645));
  OR2 U5337 ( .A(n5646), .B(n5647), .Z(n5644));
  AN2 U5338 ( .A(pi075), .B(pi156), .Z(n5647));
  AN2 U5339 ( .A(n5648), .B(n5649), .Z(n5646));
  OR2 U5340 ( .A(pi075), .B(pi156), .Z(n5649));
  OR2 U5341 ( .A(n5650), .B(n5651), .Z(n5648));
  AN2 U5342 ( .A(pi040), .B(n5652), .Z(n5651));
  AN2 U5343 ( .A(pi047), .B(n5653), .Z(n5650));
  OR2 U5344 ( .A(pi040), .B(n5652), .Z(n5653));
  AN2 U5345 ( .A(pi192), .B(n5654), .Z(n5635));
  OR2 U5346 ( .A(n5655), .B(n5656), .Z(n5654));
  OR2 U5347 ( .A(n5657), .B(n5658), .Z(n5656));
  AN2 U5348 ( .A(pi101), .B(n5659), .Z(n5658));
  AN2 U5349 ( .A(n5660), .B(n4628), .Z(n5657));
  OR2 U5350 ( .A(n5661), .B(n5659), .Z(n5660));
  OR2 U5351 ( .A(n5662), .B(n5663), .Z(n5659));
  AN2 U5352 ( .A(n5664), .B(pi036), .Z(n5663));
  AN2 U5353 ( .A(n5665), .B(n4861), .Z(n5662));
  OR2 U5354 ( .A(n5666), .B(n5664), .Z(n5665));
  AN2 U5355 ( .A(n5667), .B(n5668), .Z(n5664));
  IV2 U5356 ( .A(n5669), .Z(n5668));
  AN2 U5357 ( .A(n5670), .B(n5671), .Z(n5669));
  OR2 U5358 ( .A(po039), .B(n5672), .Z(n5671));
  AN2 U5359 ( .A(n5673), .B(n5331), .Z(n5672));
  OR2 U5360 ( .A(n5673), .B(n5331), .Z(n5670));
  IV2 U5361 ( .A(pi168), .Z(n5331));
  IV2 U5362 ( .A(n5652), .Z(n5673));
  OR2 U5363 ( .A(n5674), .B(n5675), .Z(n5652));
  AN2 U5364 ( .A(n5676), .B(n2837), .Z(n5675));
  OR2 U5365 ( .A(n5677), .B(n5678), .Z(n5676));
  AN2 U5366 ( .A(pi143), .B(pi108), .Z(n5678));
  AN2 U5367 ( .A(n5679), .B(n5680), .Z(n5677));
  OR2 U5368 ( .A(pi108), .B(pi143), .Z(n5680));
  OR2 U5369 ( .A(n5681), .B(n5682), .Z(n5679));
  AN2 U5370 ( .A(pi014), .B(pi114), .Z(n5682));
  AN2 U5371 ( .A(n5683), .B(n5684), .Z(n5681));
  OR2 U5372 ( .A(pi014), .B(pi114), .Z(n5684));
  OR2 U5373 ( .A(n5685), .B(n5686), .Z(n5683));
  OR2 U5374 ( .A(n5687), .B(n5688), .Z(n5686));
  AN2 U5375 ( .A(n5689), .B(pi170), .Z(n5688));
  AN2 U5376 ( .A(pi176), .B(n5690), .Z(n5687));
  OR2 U5377 ( .A(n5691), .B(n5689), .Z(n5690));
  AN2 U5378 ( .A(n5692), .B(n5693), .Z(n5689));
  IV2 U5379 ( .A(n5694), .Z(n5693));
  AN2 U5380 ( .A(n5695), .B(n5696), .Z(n5694));
  OR2 U5381 ( .A(n5697), .B(n4899), .Z(n5696));
  IV2 U5382 ( .A(pi097), .Z(n4899));
  AN2 U5383 ( .A(n5698), .B(n4077), .Z(n5697));
  OR2 U5384 ( .A(n5698), .B(n4077), .Z(n5695));
  AN2 U5385 ( .A(pi170), .B(n5692), .Z(n5691));
  OR2 U5386 ( .A(pi160), .B(pi189), .Z(n5692));
  AN2 U5387 ( .A(pi189), .B(pi160), .Z(n5685));
  AN2 U5388 ( .A(pi192), .B(n5699), .Z(n5674));
  OR2 U5389 ( .A(n5700), .B(n5701), .Z(n5699));
  AN2 U5390 ( .A(pi089), .B(n4881), .Z(n5701));
  AN2 U5391 ( .A(n5702), .B(n5703), .Z(n5700));
  OR2 U5392 ( .A(pi089), .B(n4881), .Z(n5703));
  OR2 U5393 ( .A(n5704), .B(n5705), .Z(n5702));
  AN2 U5394 ( .A(pi027), .B(n4885), .Z(n5705));
  AN2 U5395 ( .A(n5706), .B(n5707), .Z(n5704));
  OR2 U5396 ( .A(pi027), .B(n4885), .Z(n5707));
  OR2 U5397 ( .A(n5708), .B(n5709), .Z(n5706));
  OR2 U5398 ( .A(n5710), .B(n5711), .Z(n5709));
  AN2 U5399 ( .A(n5712), .B(pi083), .Z(n5711));
  AN2 U5400 ( .A(n5713), .B(n4877), .Z(n5710));
  OR2 U5401 ( .A(n5714), .B(n5712), .Z(n5713));
  AN2 U5402 ( .A(n5715), .B(n5716), .Z(n5712));
  IV2 U5403 ( .A(n5717), .Z(n5716));
  AN2 U5404 ( .A(n5718), .B(n5719), .Z(n5717));
  OR2 U5405 ( .A(po025), .B(n5720), .Z(n5719));
  AN2 U5406 ( .A(n5698), .B(n5303), .Z(n5720));
  OR2 U5407 ( .A(n5698), .B(n5303), .Z(n5718));
  IV2 U5408 ( .A(pi140), .Z(n5303));
  IV2 U5409 ( .A(n5721), .Z(n5698));
  OR2 U5410 ( .A(n5722), .B(n5723), .Z(n5721));
  AN2 U5411 ( .A(n5724), .B(n2837), .Z(n5723));
  OR2 U5412 ( .A(n5725), .B(n5726), .Z(n5724));
  OR2 U5413 ( .A(n5727), .B(n5728), .Z(n5726));
  AN2 U5414 ( .A(n5729), .B(pi094), .Z(n5728));
  AN2 U5415 ( .A(pi128), .B(n5730), .Z(n5727));
  OR2 U5416 ( .A(n5731), .B(n5729), .Z(n5730));
  AN2 U5417 ( .A(n5732), .B(n5733), .Z(n5729));
  IV2 U5418 ( .A(n5734), .Z(n5733));
  AN2 U5419 ( .A(n5735), .B(n5736), .Z(n5734));
  OR2 U5420 ( .A(n5737), .B(n5738), .Z(n5736));
  AN2 U5421 ( .A(n5739), .B(n5740), .Z(n5738));
  OR2 U5422 ( .A(n5741), .B(n5115), .Z(n5740));
  AN2 U5423 ( .A(n5742), .B(n4778), .Z(n5741));
  OR2 U5424 ( .A(n5742), .B(n4778), .Z(n5739));
  IV2 U5425 ( .A(pi163), .Z(n4778));
  AN2 U5426 ( .A(n3177), .B(n4770), .Z(n5737));
  OR2 U5427 ( .A(n3177), .B(n4770), .Z(n5735));
  IV2 U5428 ( .A(pi028), .Z(n4770));
  AN2 U5429 ( .A(pi094), .B(n5732), .Z(n5731));
  OR2 U5430 ( .A(pi173), .B(pi185), .Z(n5732));
  AN2 U5431 ( .A(pi173), .B(pi185), .Z(n5725));
  AN2 U5432 ( .A(pi192), .B(n5743), .Z(n5722));
  OR2 U5433 ( .A(n5744), .B(n5745), .Z(n5743));
  OR2 U5434 ( .A(n5746), .B(n5747), .Z(n5745));
  AN2 U5435 ( .A(pi131), .B(n5748), .Z(n5747));
  AN2 U5436 ( .A(n5749), .B(n5040), .Z(n5746));
  OR2 U5437 ( .A(n5750), .B(n5748), .Z(n5749));
  OR2 U5438 ( .A(n5751), .B(n5752), .Z(n5748));
  AN2 U5439 ( .A(n5753), .B(pi059), .Z(n5752));
  AN2 U5440 ( .A(n5754), .B(n3286), .Z(n5751));
  OR2 U5441 ( .A(n5755), .B(n5753), .Z(n5754));
  AN2 U5442 ( .A(n5756), .B(n5757), .Z(n5753));
  IV2 U5443 ( .A(n5758), .Z(n5757));
  AN2 U5444 ( .A(n5759), .B(n5760), .Z(n5758));
  OR2 U5445 ( .A(po010), .B(n5761), .Z(n5760));
  AN2 U5446 ( .A(n5742), .B(n5439), .Z(n5761));
  OR2 U5447 ( .A(n5742), .B(n5439), .Z(n5759));
  IV2 U5448 ( .A(pi197), .Z(n5439));
  IV2 U5449 ( .A(n5762), .Z(n5742));
  OR2 U5450 ( .A(n5763), .B(n5764), .Z(n5762));
  AN2 U5451 ( .A(n5765), .B(n2837), .Z(n5764));
  OR2 U5452 ( .A(n5766), .B(n5767), .Z(n5765));
  AN2 U5453 ( .A(pi021), .B(pi201), .Z(n5767));
  AN2 U5454 ( .A(n5768), .B(n5769), .Z(n5766));
  OR2 U5455 ( .A(pi021), .B(pi201), .Z(n5769));
  OR2 U5456 ( .A(n5770), .B(n5771), .Z(n5768));
  IV2 U5457 ( .A(n5772), .Z(n5771));
  AN2 U5458 ( .A(n5773), .B(n5774), .Z(n5772));
  OR2 U5459 ( .A(n5775), .B(n5022), .Z(n5774));
  OR2 U5460 ( .A(n5431), .B(n5776), .Z(n5773));
  AN2 U5461 ( .A(n5777), .B(n5775), .Z(n5776));
  OR2 U5462 ( .A(n5778), .B(n5779), .Z(n5775));
  AN2 U5463 ( .A(n5780), .B(n5781), .Z(n5779));
  OR2 U5464 ( .A(n5782), .B(n5783), .Z(n5781));
  AN2 U5465 ( .A(n5784), .B(n5785), .Z(n5783));
  OR2 U5466 ( .A(n5786), .B(n5787), .Z(n5785));
  IV2 U5467 ( .A(pi181), .Z(n5787));
  AN2 U5468 ( .A(n2982), .B(n5019), .Z(n5786));
  OR2 U5469 ( .A(n2982), .B(n5019), .Z(n5784));
  IV2 U5470 ( .A(pi011), .Z(n5019));
  AN2 U5471 ( .A(n5027), .B(n2957), .Z(n5782));
  OR2 U5472 ( .A(n2957), .B(n5027), .Z(n5780));
  IV2 U5473 ( .A(pi086), .Z(n5027));
  OR2 U5474 ( .A(n5022), .B(n5778), .Z(n5777));
  AN2 U5475 ( .A(n5165), .B(n5031), .Z(n5778));
  IV2 U5476 ( .A(pi165), .Z(n5031));
  IV2 U5477 ( .A(pi032), .Z(n5022));
  AN2 U5478 ( .A(pi165), .B(pi107), .Z(n5770));
  AN2 U5479 ( .A(pi192), .B(n5788), .Z(n5763));
  OR2 U5480 ( .A(n5789), .B(n5790), .Z(n5788));
  AN2 U5481 ( .A(pi121), .B(n5000), .Z(n5790));
  AN2 U5482 ( .A(n5791), .B(n5792), .Z(n5789));
  OR2 U5483 ( .A(pi121), .B(n5000), .Z(n5792));
  OR2 U5484 ( .A(n5793), .B(n5794), .Z(n5791));
  AN2 U5485 ( .A(pi053), .B(n5795), .Z(n5794));
  AN2 U5486 ( .A(n5796), .B(n5004), .Z(n5793));
  OR2 U5487 ( .A(pi053), .B(n5795), .Z(n5796));
  OR2 U5488 ( .A(n5797), .B(n5798), .Z(n5795));
  AN2 U5489 ( .A(pi184), .B(n5008), .Z(n5798));
  AN2 U5490 ( .A(n5799), .B(n5800), .Z(n5797));
  OR2 U5491 ( .A(pi184), .B(n5008), .Z(n5800));
  OR2 U5492 ( .A(n5801), .B(n5802), .Z(n5799));
  AN2 U5493 ( .A(pi181), .B(pi103), .Z(n5802));
  AN2 U5494 ( .A(n5803), .B(n2962), .Z(n5801));
  OR2 U5495 ( .A(pi103), .B(pi181), .Z(n5803));
  AN2 U5496 ( .A(pi059), .B(n5756), .Z(n5755));
  AN2 U5497 ( .A(pi131), .B(n5756), .Z(n5750));
  OR2 U5498 ( .A(pi001), .B(n5037), .Z(n5756));
  AN2 U5499 ( .A(pi001), .B(n5037), .Z(n5744));
  AN2 U5500 ( .A(pi083), .B(n5715), .Z(n5714));
  OR2 U5501 ( .A(pi162), .B(n4874), .Z(n5715));
  AN2 U5502 ( .A(pi162), .B(n4874), .Z(n5708));
  AN2 U5503 ( .A(pi036), .B(n5667), .Z(n5666));
  AN2 U5504 ( .A(pi101), .B(n5667), .Z(n5661));
  OR2 U5505 ( .A(pi205), .B(n4915), .Z(n5667));
  AN2 U5506 ( .A(pi205), .B(n4915), .Z(n5655));
  AN2 U5507 ( .A(po036), .B(n5350), .Z(n5630));
  OR2 U5508 ( .A(po036), .B(n5350), .Z(n5628));
  IV2 U5509 ( .A(pi018), .Z(n5350));
  AN2 U5510 ( .A(pi099), .B(n5625), .Z(n5624));
  OR2 U5511 ( .A(pi180), .B(n4947), .Z(n5625));
  AN2 U5512 ( .A(pi180), .B(n4947), .Z(n5618));
  AN2 U5513 ( .A(n3261), .B(pi049), .Z(n5347));
  AN2 U5514 ( .A(n3926), .B(n5804), .Z(n5551));
  OR2 U5515 ( .A(n5805), .B(n5806), .Z(n5804));
  OR2 U5516 ( .A(pi085), .B(pi019), .Z(n5806));
  OR2 U5517 ( .A(pi110), .B(n5807), .Z(n5805));
  OR2 U5518 ( .A(pi167), .B(pi164), .Z(n5807));
  AN2 U5519 ( .A(pi126), .B(pi190), .Z(n5549));
  AN2 U5520 ( .A(n5808), .B(pi035), .Z(n5547));
  AN2 U5521 ( .A(pi056), .B(pi100), .Z(n5808));
  AN2 U5522 ( .A(pi054), .B(n5809), .Z(n5504));
  OR2 U5523 ( .A(n4167), .B(n5810), .Z(n5809));
  OR2 U5524 ( .A(pi146), .B(pi025), .Z(n5810));
  AN2 U5525 ( .A(n5811), .B(n2882), .Z(po017));
  OR2 U5526 ( .A(pi200), .B(n3003), .Z(n5811));
  OR2 U5527 ( .A(n5812), .B(n5813), .Z(po016));
  OR2 U5528 ( .A(n5814), .B(n5815), .Z(n5813));
  AN2 U5529 ( .A(n3280), .B(n3064), .Z(n5815));
  AN2 U5530 ( .A(n5100), .B(n5816), .Z(n5814));
  OR2 U5531 ( .A(n5817), .B(n5818), .Z(n5816));
  AN2 U5532 ( .A(n3055), .B(n5819), .Z(n5818));
  OR2 U5533 ( .A(n2845), .B(n3143), .Z(n5819));
  OR2 U5534 ( .A(n2978), .B(n3147), .Z(n3143));
  AN2 U5535 ( .A(n3127), .B(n5820), .Z(n5817));
  OR2 U5536 ( .A(n2833), .B(n3138), .Z(n5820));
  OR2 U5537 ( .A(n2880), .B(n3147), .Z(n3138));
  OR2 U5538 ( .A(n2998), .B(n5821), .Z(n3147));
  OR2 U5539 ( .A(n2882), .B(n2862), .Z(n5821));
  OR2 U5540 ( .A(n2925), .B(n2901), .Z(n2882));
  AN2 U5541 ( .A(pi192), .B(n3036), .Z(n3127));
  IV2 U5542 ( .A(n5822), .Z(n5100));
  OR2 U5543 ( .A(n5823), .B(n5824), .Z(n5812));
  AN2 U5544 ( .A(n5825), .B(pi192), .Z(n5824));
  AN2 U5545 ( .A(n5826), .B(po010), .Z(n5825));
  AN2 U5546 ( .A(n5827), .B(n2837), .Z(n5823));
  AN2 U5547 ( .A(n5828), .B(n5829), .Z(n5827));
  OR2 U5548 ( .A(n5830), .B(n5831), .Z(po008));
  AN2 U5549 ( .A(n3344), .B(n3251), .Z(n5831));
  OR2 U5550 ( .A(n5832), .B(n5833), .Z(n3251));
  AN2 U5551 ( .A(n3355), .B(n5454), .Z(n5832));
  OR2 U5552 ( .A(n5834), .B(n5835), .Z(n5454));
  AN2 U5553 ( .A(n5836), .B(n4426), .Z(n5834));
  IV2 U5554 ( .A(n3352), .Z(n3355));
  AN2 U5555 ( .A(n3250), .B(n5837), .Z(n5830));
  OR2 U5556 ( .A(n5838), .B(n5839), .Z(n5837));
  OR2 U5557 ( .A(n5840), .B(n3245), .Z(n5839));
  OR2 U5558 ( .A(n5841), .B(n5842), .Z(n3245));
  AN2 U5559 ( .A(n3244), .B(n3699), .Z(n5842));
  AN2 U5560 ( .A(n3242), .B(n3700), .Z(n5841));
  IV2 U5561 ( .A(n5843), .Z(n3242));
  AN2 U5562 ( .A(n3352), .B(n3701), .Z(n5840));
  OR2 U5563 ( .A(n5844), .B(n5845), .Z(n5838));
  AN2 U5564 ( .A(n4418), .B(n3762), .Z(n5845));
  AN2 U5565 ( .A(n5846), .B(n3236), .Z(n5844));
  OR2 U5566 ( .A(pi037), .B(n5847), .Z(po007));
  IV2 U5567 ( .A(pi116), .Z(n5847));
  OR2 U5568 ( .A(n5848), .B(n5849), .Z(po006));
  AN2 U5569 ( .A(n3370), .B(n5850), .Z(n5849));
  OR2 U5570 ( .A(n5851), .B(n5852), .Z(n5850));
  OR2 U5571 ( .A(n5853), .B(n5138), .Z(n5852));
  OR2 U5572 ( .A(n5854), .B(n3566), .Z(n5138));
  AN2 U5573 ( .A(n3512), .B(n3926), .Z(n3566));
  AN2 U5574 ( .A(n3926), .B(n4368), .Z(n5854));
  OR2 U5575 ( .A(n5855), .B(n5856), .Z(n5851));
  AN2 U5576 ( .A(n5139), .B(n3380), .Z(n5856));
  OR2 U5577 ( .A(n5857), .B(n5858), .Z(n5139));
  AN2 U5578 ( .A(n5859), .B(n3261), .Z(n5857));
  AN2 U5579 ( .A(n5860), .B(pi118), .Z(n5855));
  AN2 U5580 ( .A(n5861), .B(n3261), .Z(n5860));
  OR2 U5581 ( .A(n5858), .B(n5859), .Z(n5861));
  OR2 U5582 ( .A(n5862), .B(n5863), .Z(n5859));
  OR2 U5583 ( .A(n3404), .B(n5864), .Z(n5863));
  AN2 U5584 ( .A(n5865), .B(pi060), .Z(n5864));
  AN2 U5585 ( .A(n4368), .B(n5866), .Z(n5865));
  IV2 U5586 ( .A(n3446), .Z(n3404));
  AN2 U5587 ( .A(n4367), .B(pi196), .Z(n5862));
  IV2 U5588 ( .A(n4364), .Z(n4367));
  IV2 U5589 ( .A(n5867), .Z(n5858));
  IV2 U5590 ( .A(n3393), .Z(n3370));
  AN2 U5591 ( .A(n3393), .B(n5868), .Z(n5848));
  OR2 U5592 ( .A(n5869), .B(n5870), .Z(n5868));
  OR2 U5593 ( .A(n5135), .B(n5871), .Z(n5870));
  AN2 U5594 ( .A(n3480), .B(n5872), .Z(n5871));
  AN2 U5595 ( .A(n5867), .B(n3321), .Z(n5135));
  OR2 U5596 ( .A(po104), .B(n4364), .Z(n5867));
  OR2 U5597 ( .A(n5873), .B(n5874), .Z(n5869));
  OR2 U5598 ( .A(n5875), .B(n5876), .Z(n5874));
  AN2 U5599 ( .A(n5877), .B(po071), .Z(n5876));
  OR2 U5600 ( .A(n5136), .B(n5878), .Z(n5877));
  OR2 U5601 ( .A(n5879), .B(n5880), .Z(n5136));
  OR2 U5602 ( .A(n5881), .B(n5882), .Z(n5880));
  AN2 U5603 ( .A(n3398), .B(n4364), .Z(n5882));
  AN2 U5604 ( .A(n4363), .B(n3419), .Z(n5879));
  AN2 U5605 ( .A(n5883), .B(n3398), .Z(n5875));
  AN2 U5606 ( .A(n3446), .B(n3533), .Z(n3398));
  AN2 U5607 ( .A(n4364), .B(n3913), .Z(n5883));
  OR2 U5608 ( .A(n4062), .B(po027), .Z(n4364));
  IV2 U5609 ( .A(n4061), .Z(n4062));
  AN2 U5610 ( .A(n3416), .B(n4363), .Z(n5873));
  IV2 U5611 ( .A(n4368), .Z(n4363));
  OR2 U5612 ( .A(n3363), .B(n4061), .Z(n4368));
  OR2 U5613 ( .A(n5884), .B(n5885), .Z(n4061));
  OR2 U5614 ( .A(n5886), .B(n5887), .Z(n5885));
  AN2 U5615 ( .A(n5888), .B(n4943), .Z(n5887));
  AN2 U5616 ( .A(n5889), .B(n3989), .Z(n5886));
  OR2 U5617 ( .A(n5890), .B(n5891), .Z(n5884));
  OR2 U5618 ( .A(n5892), .B(n3490), .Z(n5891));
  AN2 U5619 ( .A(n5893), .B(n5894), .Z(n5890));
  AN2 U5620 ( .A(n3495), .B(n5895), .Z(n5893));
  AN2 U5621 ( .A(n3446), .B(n3480), .Z(n3416));
  OR2 U5622 ( .A(po104), .B(n3942), .Z(n3446));
  OR2 U5623 ( .A(n5896), .B(n3253), .Z(po012));
  AN2 U5624 ( .A(n5897), .B(pi054), .Z(n3253));
  OR2 U5625 ( .A(n4133), .B(n5898), .Z(n5897));
  AN2 U5626 ( .A(n4127), .B(n3255), .Z(n5896));
  OR2 U5627 ( .A(pi054), .B(n5120), .Z(n3255));
  OR2 U5628 ( .A(n5899), .B(n4167), .Z(n5120));
  AN2 U5629 ( .A(n4133), .B(n4128), .Z(n5899));
  IV2 U5630 ( .A(po064), .Z(n4133));
  OR2 U5631 ( .A(n5900), .B(n4372), .Z(n4127));
  OR2 U5632 ( .A(n5901), .B(n5902), .Z(n4372));
  AN2 U5633 ( .A(n4380), .B(n4319), .Z(n5901));
  AN2 U5634 ( .A(n5903), .B(n4374), .Z(n5900));
  OR2 U5635 ( .A(n5904), .B(n5905), .Z(n4374));
  AN2 U5636 ( .A(n5906), .B(n3261), .Z(n5905));
  OR2 U5637 ( .A(n5907), .B(n5908), .Z(n5906));
  OR2 U5638 ( .A(n5909), .B(n5910), .Z(n5908));
  AN2 U5639 ( .A(n5911), .B(po103), .Z(n5910));
  AN2 U5640 ( .A(n5912), .B(pi058), .Z(n5911));
  AN2 U5641 ( .A(n5913), .B(n5914), .Z(n5912));
  AN2 U5642 ( .A(n5915), .B(n5916), .Z(n5913));
  OR2 U5643 ( .A(pi204), .B(n5917), .Z(n5916));
  AN2 U5644 ( .A(n4057), .B(n4013), .Z(n5917));
  OR2 U5645 ( .A(n5918), .B(n5919), .Z(n5915));
  AN2 U5646 ( .A(po040), .B(n3966), .Z(n5918));
  AN2 U5647 ( .A(n5920), .B(n3265), .Z(n5909));
  AN2 U5648 ( .A(n5921), .B(n5922), .Z(n5920));
  AN2 U5649 ( .A(n4057), .B(n4316), .Z(n5922));
  AN2 U5650 ( .A(n4157), .B(n5914), .Z(n5921));
  OR2 U5651 ( .A(n5923), .B(n4319), .Z(n5914));
  AN2 U5652 ( .A(pi065), .B(pi192), .Z(n5923));
  OR2 U5653 ( .A(pi204), .B(n4013), .Z(n4157));
  AN2 U5654 ( .A(n5924), .B(n4046), .Z(n5907));
  AN2 U5655 ( .A(po040), .B(n3263), .Z(n5924));
  OR2 U5656 ( .A(n5925), .B(n2837), .Z(n3263));
  AN2 U5657 ( .A(n3264), .B(pi058), .Z(n5925));
  AN2 U5658 ( .A(n4391), .B(n4319), .Z(n5904));
  AN2 U5659 ( .A(n3265), .B(n4013), .Z(n4391));
  IV2 U5660 ( .A(n4158), .Z(n5903));
  OR2 U5661 ( .A(n4312), .B(n5926), .Z(n4158));
  OR2 U5662 ( .A(n4040), .B(n4229), .Z(n5926));
  IV2 U5663 ( .A(n4184), .Z(n4229));
  OR2 U5664 ( .A(n5927), .B(n5928), .Z(n4184));
  OR2 U5665 ( .A(n5929), .B(n5930), .Z(n5928));
  AN2 U5666 ( .A(n5931), .B(n5932), .Z(n5929));
  OR2 U5667 ( .A(n5933), .B(n5934), .Z(n5932));
  AN2 U5668 ( .A(n3457), .B(n3493), .Z(n5934));
  IV2 U5669 ( .A(n3661), .Z(n3493));
  OR2 U5670 ( .A(n5935), .B(n5936), .Z(n3661));
  OR2 U5671 ( .A(n3229), .B(n3235), .Z(n5936));
  OR2 U5672 ( .A(n5937), .B(n5938), .Z(n3235));
  OR2 U5673 ( .A(n5939), .B(n5940), .Z(n5938));
  AN2 U5674 ( .A(n5452), .B(n3241), .Z(n5940));
  AN2 U5675 ( .A(n5453), .B(n3243), .Z(n5939));
  AN2 U5676 ( .A(po082), .B(n5846), .Z(n5937));
  OR2 U5677 ( .A(n5941), .B(n5942), .Z(n5846));
  AN2 U5678 ( .A(n5452), .B(n3700), .Z(n5942));
  AN2 U5679 ( .A(n3638), .B(n3635), .Z(n5452));
  IV2 U5680 ( .A(pi098), .Z(n3638));
  AN2 U5681 ( .A(n5453), .B(n3699), .Z(n5941));
  AN2 U5682 ( .A(n3597), .B(n3593), .Z(n5453));
  OR2 U5683 ( .A(n5943), .B(n5944), .Z(n3229));
  AN2 U5684 ( .A(po082), .B(n3344), .Z(n5944));
  AN2 U5685 ( .A(n3352), .B(n5945), .Z(n5943));
  OR2 U5686 ( .A(n5946), .B(n5947), .Z(n5945));
  OR2 U5687 ( .A(n3241), .B(n3243), .Z(n5947));
  AN2 U5688 ( .A(po082), .B(n3701), .Z(n5946));
  IV2 U5689 ( .A(n5833), .Z(n3701));
  OR2 U5690 ( .A(n3233), .B(n5948), .Z(n5935));
  AN2 U5691 ( .A(n3339), .B(n5949), .Z(n5948));
  AN2 U5692 ( .A(n5949), .B(po011), .Z(n3233));
  OR2 U5693 ( .A(n5950), .B(n5951), .Z(n5949));
  OR2 U5694 ( .A(n5952), .B(n5953), .Z(n5951));
  AN2 U5695 ( .A(n3241), .B(n3635), .Z(n5953));
  AN2 U5696 ( .A(n3992), .B(n3700), .Z(n3241));
  AN2 U5697 ( .A(n3632), .B(pi192), .Z(n3700));
  IV2 U5698 ( .A(pi004), .Z(n3992));
  AN2 U5699 ( .A(n3243), .B(n3593), .Z(n5952));
  OR2 U5700 ( .A(po036), .B(n4440), .Z(n3593));
  AN2 U5701 ( .A(n5372), .B(n3699), .Z(n3243));
  AN2 U5702 ( .A(po082), .B(n3762), .Z(n5950));
  OR2 U5703 ( .A(n5954), .B(n5955), .Z(n3762));
  OR2 U5704 ( .A(n5956), .B(n5957), .Z(n5955));
  AN2 U5705 ( .A(po036), .B(n5958), .Z(n5957));
  OR2 U5706 ( .A(n5959), .B(po001), .Z(n5958));
  AN2 U5707 ( .A(pi192), .B(n5960), .Z(n5956));
  OR2 U5708 ( .A(n5961), .B(n5962), .Z(n5960));
  AN2 U5709 ( .A(po001), .B(n4001), .Z(n5962));
  AN2 U5710 ( .A(n3635), .B(n3998), .Z(n5961));
  OR2 U5711 ( .A(po036), .B(n4001), .Z(n3635));
  IV2 U5712 ( .A(pi171), .Z(n4001));
  AN2 U5713 ( .A(n3699), .B(n4440), .Z(n5954));
  AN2 U5714 ( .A(n2837), .B(n3590), .Z(n3699));
  AN2 U5715 ( .A(n5963), .B(n3667), .Z(n5933));
  AN2 U5716 ( .A(n3291), .B(n3341), .Z(n3667));
  IV2 U5717 ( .A(n3339), .Z(n3341));
  OR2 U5718 ( .A(n5964), .B(n5965), .Z(n3339));
  AN2 U5719 ( .A(n5966), .B(n4441), .Z(n5965));
  AN2 U5720 ( .A(n5448), .B(po036), .Z(n5964));
  IV2 U5721 ( .A(n5966), .Z(n5448));
  OR2 U5722 ( .A(n5967), .B(n5968), .Z(n3291));
  AN2 U5723 ( .A(n5969), .B(n3688), .Z(n5968));
  IV2 U5724 ( .A(n3746), .Z(n5969));
  AN2 U5725 ( .A(po011), .B(n3746), .Z(n5967));
  OR2 U5726 ( .A(n3717), .B(n3705), .Z(n3746));
  AN2 U5727 ( .A(n3495), .B(n5970), .Z(n5963));
  OR2 U5728 ( .A(n5971), .B(n5972), .Z(n5970));
  OR2 U5729 ( .A(n5973), .B(n5974), .Z(n5972));
  AN2 U5730 ( .A(n5975), .B(pi192), .Z(n5974));
  AN2 U5731 ( .A(n3567), .B(n5976), .Z(n5975));
  OR2 U5732 ( .A(n5977), .B(n5978), .Z(n5976));
  OR2 U5733 ( .A(n5979), .B(n5980), .Z(n5978));
  AN2 U5734 ( .A(n4635), .B(n5981), .Z(n5979));
  IV2 U5735 ( .A(n4464), .Z(n4635));
  OR2 U5736 ( .A(po039), .B(n3870), .Z(n4464));
  IV2 U5737 ( .A(pi016), .Z(n3870));
  OR2 U5738 ( .A(n5982), .B(n5983), .Z(n5977));
  AN2 U5739 ( .A(n5984), .B(n3033), .Z(n5983));
  IV2 U5740 ( .A(n3038), .Z(n3033));
  OR2 U5741 ( .A(po070), .B(n3199), .Z(n3038));
  IV2 U5742 ( .A(pi096), .Z(n3199));
  AN2 U5743 ( .A(n5985), .B(n5986), .Z(n5982));
  OR2 U5744 ( .A(n5987), .B(n3042), .Z(n5986));
  IV2 U5745 ( .A(n3037), .Z(n3042));
  OR2 U5746 ( .A(po099), .B(n3171), .Z(n3037));
  AN2 U5747 ( .A(n3063), .B(n5988), .Z(n5987));
  OR2 U5748 ( .A(n5989), .B(n5990), .Z(n5988));
  AN2 U5749 ( .A(n3036), .B(n5991), .Z(n5989));
  OR2 U5750 ( .A(n5992), .B(n3010), .Z(n5991));
  OR2 U5751 ( .A(n5993), .B(n5994), .Z(n3010));
  AN2 U5752 ( .A(pi088), .B(n3012), .Z(n5992));
  IV2 U5753 ( .A(n5995), .Z(n3036));
  OR2 U5754 ( .A(n5996), .B(n5990), .Z(n5995));
  AN2 U5755 ( .A(pi166), .B(n3049), .Z(n5990));
  AN2 U5756 ( .A(po010), .B(n3106), .Z(n5996));
  OR2 U5757 ( .A(n3534), .B(n3363), .Z(n3567));
  AN2 U5758 ( .A(n5997), .B(n3457), .Z(n5973));
  IV2 U5759 ( .A(n4060), .Z(n3457));
  OR2 U5760 ( .A(n5998), .B(n5999), .Z(n4060));
  AN2 U5761 ( .A(po027), .B(n3451), .Z(n5998));
  AN2 U5762 ( .A(n3760), .B(n4652), .Z(n5997));
  AN2 U5763 ( .A(n6000), .B(n6001), .Z(n5971));
  OR2 U5764 ( .A(n3261), .B(n3525), .Z(n6001));
  AN2 U5765 ( .A(n3363), .B(n3321), .Z(n3525));
  OR2 U5766 ( .A(n6002), .B(n6003), .Z(n6000));
  AN2 U5767 ( .A(n6004), .B(n2837), .Z(n6003));
  OR2 U5768 ( .A(n6005), .B(n6006), .Z(n6004));
  OR2 U5769 ( .A(n6007), .B(n6008), .Z(n6006));
  AN2 U5770 ( .A(n4641), .B(n5981), .Z(n6007));
  IV2 U5771 ( .A(n4468), .Z(n4641));
  OR2 U5772 ( .A(po039), .B(n4735), .Z(n4468));
  IV2 U5773 ( .A(pi040), .Z(n4735));
  OR2 U5774 ( .A(n6009), .B(n6010), .Z(n6005));
  AN2 U5775 ( .A(n5985), .B(n6011), .Z(n6010));
  OR2 U5776 ( .A(n6012), .B(n6013), .Z(n6011));
  OR2 U5777 ( .A(n3066), .B(n6014), .Z(n6013));
  AN2 U5778 ( .A(n6015), .B(n6016), .Z(n6014));
  IV2 U5779 ( .A(n3112), .Z(n3066));
  OR2 U5780 ( .A(po099), .B(n3177), .Z(n3112));
  AN2 U5781 ( .A(n6017), .B(n6018), .Z(n6012));
  OR2 U5782 ( .A(n6019), .B(n6020), .Z(n6018));
  AN2 U5783 ( .A(n6021), .B(n3119), .Z(n6019));
  OR2 U5784 ( .A(n6022), .B(n5993), .Z(n6021));
  AN2 U5785 ( .A(n2890), .B(n5000), .Z(n5993));
  AN2 U5786 ( .A(pi201), .B(n3012), .Z(n6022));
  OR2 U5787 ( .A(n2890), .B(n5000), .Z(n3012));
  IV2 U5788 ( .A(n2886), .Z(n2890));
  OR2 U5789 ( .A(n6023), .B(n6024), .Z(n2886));
  OR2 U5790 ( .A(n6025), .B(n6026), .Z(n6024));
  AN2 U5791 ( .A(n6027), .B(n2998), .Z(n6026));
  AN2 U5792 ( .A(po079), .B(n6028), .Z(n6025));
  OR2 U5793 ( .A(n6029), .B(n4095), .Z(n6028));
  OR2 U5794 ( .A(n6030), .B(n6031), .Z(n4095));
  AN2 U5795 ( .A(n4098), .B(n2887), .Z(n6031));
  AN2 U5796 ( .A(n6032), .B(po031), .Z(n6030));
  AN2 U5797 ( .A(n2990), .B(n2974), .Z(n6032));
  AN2 U5798 ( .A(n2990), .B(n5169), .Z(n6029));
  OR2 U5799 ( .A(n6033), .B(po106), .Z(n2990));
  AN2 U5800 ( .A(n2837), .B(n5431), .Z(n6033));
  OR2 U5801 ( .A(n6034), .B(n6035), .Z(n6023));
  AN2 U5802 ( .A(n4099), .B(n6036), .Z(n6035));
  OR2 U5803 ( .A(n6037), .B(n6038), .Z(n6036));
  AN2 U5804 ( .A(n6039), .B(n5165), .Z(n6038));
  OR2 U5805 ( .A(n6040), .B(n5169), .Z(n6039));
  OR2 U5806 ( .A(n2978), .B(n2862), .Z(n5169));
  AN2 U5807 ( .A(po031), .B(n2974), .Z(n6040));
  AN2 U5808 ( .A(n6041), .B(n2974), .Z(n6037));
  AN2 U5809 ( .A(n5172), .B(n2957), .Z(n6041));
  AN2 U5810 ( .A(n2947), .B(n2837), .Z(n4099));
  AN2 U5811 ( .A(n6042), .B(n4098), .Z(n6034));
  AN2 U5812 ( .A(n2891), .B(pi192), .Z(n4098));
  IV2 U5813 ( .A(n2892), .Z(n2891));
  AN2 U5814 ( .A(n6043), .B(n3847), .Z(n6042));
  IV2 U5815 ( .A(n2885), .Z(n6043));
  AN2 U5816 ( .A(n5984), .B(n3076), .Z(n6009));
  IV2 U5817 ( .A(n3109), .Z(n3076));
  OR2 U5818 ( .A(po070), .B(n3205), .Z(n3109));
  IV2 U5819 ( .A(pi128), .Z(n3205));
  AN2 U5820 ( .A(n5985), .B(n6044), .Z(n6002));
  OR2 U5821 ( .A(n6045), .B(n6046), .Z(n5927));
  AN2 U5822 ( .A(n6047), .B(n3945), .Z(n6046));
  IV2 U5823 ( .A(n4313), .Z(n3945));
  OR2 U5824 ( .A(n3321), .B(n2837), .Z(n4313));
  AN2 U5825 ( .A(pi050), .B(n4975), .Z(n6047));
  AN2 U5826 ( .A(n6048), .B(n6049), .Z(n6045));
  AN2 U5827 ( .A(n6050), .B(n6051), .Z(n6049));
  OR2 U5828 ( .A(n3363), .B(n6052), .Z(n6051));
  OR2 U5829 ( .A(po027), .B(n3989), .Z(n6050));
  AN2 U5830 ( .A(n6053), .B(n4943), .Z(n6048));
  OR2 U5831 ( .A(n4239), .B(n4192), .Z(n4312));
  OR2 U5832 ( .A(n6054), .B(n6055), .Z(po003));
  OR2 U5833 ( .A(n6056), .B(n6057), .Z(n6055));
  AN2 U5834 ( .A(n6058), .B(pi054), .Z(n6057));
  OR2 U5835 ( .A(n6059), .B(n6060), .Z(n6058));
  AN2 U5836 ( .A(n4177), .B(n5126), .Z(n6060));
  AN2 U5837 ( .A(n5125), .B(n5898), .Z(n6059));
  AN2 U5838 ( .A(n6061), .B(n4129), .Z(n6056));
  AN2 U5839 ( .A(n4177), .B(n5125), .Z(n6061));
  OR2 U5840 ( .A(n6062), .B(n3257), .Z(n5125));
  OR2 U5841 ( .A(n5902), .B(n6063), .Z(n3257));
  OR2 U5842 ( .A(n6064), .B(n6065), .Z(n6063));
  AN2 U5843 ( .A(n4403), .B(n4319), .Z(n6065));
  IV2 U5844 ( .A(po004), .Z(n4319));
  OR2 U5845 ( .A(n6066), .B(n4380), .Z(n4403));
  AN2 U5846 ( .A(n6067), .B(n3259), .Z(n6066));
  AN2 U5847 ( .A(n4053), .B(n4013), .Z(n6067));
  OR2 U5848 ( .A(n6068), .B(n3265), .Z(n4053));
  AN2 U5849 ( .A(pi058), .B(n3261), .Z(n6068));
  AN2 U5850 ( .A(n6069), .B(n6070), .Z(n6064));
  AN2 U5851 ( .A(n4387), .B(n4013), .Z(n6070));
  IV2 U5852 ( .A(po040), .Z(n4013));
  AN2 U5853 ( .A(pi065), .B(n3259), .Z(n6069));
  OR2 U5854 ( .A(n6071), .B(n4379), .Z(n5902));
  IV2 U5855 ( .A(n4159), .Z(n4379));
  AN2 U5856 ( .A(n4380), .B(n4404), .Z(n6071));
  IV2 U5857 ( .A(n4161), .Z(n4404));
  IV2 U5858 ( .A(n4141), .Z(n4380));
  OR2 U5859 ( .A(n4016), .B(n6072), .Z(n4141));
  OR2 U5860 ( .A(n6073), .B(n6074), .Z(n6072));
  AN2 U5861 ( .A(n6075), .B(n4242), .Z(n6074));
  OR2 U5862 ( .A(n6076), .B(n6077), .Z(n4016));
  AN2 U5863 ( .A(n4040), .B(n3951), .Z(n6076));
  AN2 U5864 ( .A(n3259), .B(n6078), .Z(n6062));
  OR2 U5865 ( .A(n6079), .B(n3926), .Z(n6078));
  AN2 U5866 ( .A(n3264), .B(n4387), .Z(n6079));
  AN2 U5867 ( .A(n3261), .B(n4026), .Z(n4387));
  IV2 U5868 ( .A(n6080), .Z(n3264));
  OR2 U5869 ( .A(n6081), .B(n5919), .Z(n6080));
  AN2 U5870 ( .A(n4330), .B(n6082), .Z(n3259));
  AN2 U5871 ( .A(n4205), .B(n3314), .Z(n6082));
  IV2 U5872 ( .A(n5898), .Z(n4177));
  AN2 U5873 ( .A(n4172), .B(n5126), .Z(n6054));
  OR2 U5874 ( .A(n6083), .B(n6084), .Z(n5126));
  OR2 U5875 ( .A(n6085), .B(n6086), .Z(n6084));
  AN2 U5876 ( .A(n4227), .B(n4159), .Z(n6086));
  OR2 U5877 ( .A(po004), .B(n4161), .Z(n4159));
  OR2 U5878 ( .A(n4310), .B(n3321), .Z(n4161));
  OR2 U5879 ( .A(n6087), .B(n6088), .Z(n4227));
  OR2 U5880 ( .A(n6089), .B(n6077), .Z(n6088));
  OR2 U5881 ( .A(n6090), .B(n6091), .Z(n6077));
  OR2 U5882 ( .A(n3317), .B(n6092), .Z(n6091));
  AN2 U5883 ( .A(n4291), .B(n4056), .Z(n6092));
  AN2 U5884 ( .A(n3321), .B(po103), .Z(n3317));
  AN2 U5885 ( .A(n4040), .B(n3321), .Z(n6090));
  AN2 U5886 ( .A(n4192), .B(n6075), .Z(n6089));
  OR2 U5887 ( .A(n3321), .B(n6093), .Z(n6075));
  OR2 U5888 ( .A(n6073), .B(n6094), .Z(n6087));
  AN2 U5889 ( .A(n4040), .B(n4291), .Z(n6094));
  AN2 U5890 ( .A(po040), .B(n6095), .Z(n6073));
  OR2 U5891 ( .A(n4040), .B(n6096), .Z(n6095));
  OR2 U5892 ( .A(n3318), .B(n4293), .Z(n6096));
  OR2 U5893 ( .A(n3951), .B(n3321), .Z(n4293));
  AN2 U5894 ( .A(n4056), .B(n6097), .Z(n3318));
  AN2 U5895 ( .A(n4057), .B(pi192), .Z(n6097));
  IV2 U5896 ( .A(n4026), .Z(n4056));
  OR2 U5897 ( .A(pi058), .B(n3265), .Z(n4026));
  IV2 U5898 ( .A(n3314), .Z(n4040));
  OR2 U5899 ( .A(n6098), .B(n4201), .Z(n3314));
  IV2 U5900 ( .A(po091), .Z(n4201));
  AN2 U5901 ( .A(n3261), .B(n4200), .Z(n6098));
  AN2 U5902 ( .A(n6081), .B(pi192), .Z(n6085));
  AN2 U5903 ( .A(n4150), .B(po004), .Z(n6081));
  IV2 U5904 ( .A(pi065), .Z(n4150));
  OR2 U5905 ( .A(n6099), .B(n4396), .Z(n6083));
  AN2 U5906 ( .A(n4406), .B(n6100), .Z(n4396));
  OR2 U5907 ( .A(n6101), .B(n3321), .Z(n6100));
  AN2 U5908 ( .A(n6102), .B(n6103), .Z(n6101));
  AN2 U5909 ( .A(n4223), .B(n4057), .Z(n6103));
  AN2 U5910 ( .A(n4310), .B(n6104), .Z(n6102));
  OR2 U5911 ( .A(po040), .B(n5919), .Z(n6104));
  IV2 U5912 ( .A(pi204), .Z(n5919));
  IV2 U5913 ( .A(n4156), .Z(n4310));
  OR2 U5914 ( .A(pi065), .B(n2837), .Z(n4156));
  AN2 U5915 ( .A(po004), .B(n6105), .Z(n6099));
  OR2 U5916 ( .A(n6106), .B(n3321), .Z(n6105));
  AN2 U5917 ( .A(n4406), .B(n6093), .Z(n6106));
  OR2 U5918 ( .A(n6107), .B(n4028), .Z(n6093));
  AN2 U5919 ( .A(n4223), .B(n4291), .Z(n4028));
  AN2 U5920 ( .A(n4057), .B(n3951), .Z(n4291));
  IV2 U5921 ( .A(n4041), .Z(n3951));
  OR2 U5922 ( .A(pi204), .B(n2837), .Z(n4041));
  OR2 U5923 ( .A(po103), .B(n4316), .Z(n4223));
  IV2 U5924 ( .A(pi058), .Z(n4316));
  AN2 U5925 ( .A(po040), .B(n3322), .Z(n6107));
  OR2 U5926 ( .A(n4046), .B(n4045), .Z(n3322));
  OR2 U5927 ( .A(n6108), .B(n6109), .Z(n4045));
  AN2 U5928 ( .A(n4148), .B(n4057), .Z(n6109));
  OR2 U5929 ( .A(po091), .B(n3966), .Z(n4057));
  IV2 U5930 ( .A(pi129), .Z(n3966));
  AN2 U5931 ( .A(n4203), .B(po103), .Z(n6108));
  IV2 U5932 ( .A(n4200), .Z(n4203));
  OR2 U5933 ( .A(pi129), .B(n2837), .Z(n4200));
  AN2 U5934 ( .A(po103), .B(po091), .Z(n4046));
  AN2 U5935 ( .A(n5898), .B(n4129), .Z(n4172));
  IV2 U5936 ( .A(pi054), .Z(n4129));
  OR2 U5937 ( .A(n4167), .B(n4128), .Z(n5898));
  IV2 U5938 ( .A(po085), .Z(n4128));
  IV2 U5939 ( .A(pi052), .Z(n4167));
  AN2 U5940 ( .A(n6110), .B(n6111), .Z(po002));
  OR2 U5941 ( .A(n3306), .B(n4450), .Z(n6111));
  OR2 U5942 ( .A(n4458), .B(n4606), .Z(n6110));
  IV2 U5943 ( .A(n3306), .Z(n4458));
  OR2 U5944 ( .A(n6112), .B(n4652), .Z(n3306));
  OR2 U5945 ( .A(n6113), .B(n6114), .Z(n4652));
  AN2 U5946 ( .A(n6115), .B(n2837), .Z(n6114));
  OR2 U5947 ( .A(n6116), .B(n6117), .Z(n6115));
  AN2 U5948 ( .A(pi108), .B(n4881), .Z(n6117));
  AN2 U5949 ( .A(n4475), .B(n6118), .Z(n6116));
  OR2 U5950 ( .A(n5467), .B(n6119), .Z(n6118));
  IV2 U5951 ( .A(n5488), .Z(n6119));
  OR2 U5952 ( .A(po102), .B(n5322), .Z(n5488));
  IV2 U5953 ( .A(pi114), .Z(n5322));
  AN2 U5954 ( .A(n6120), .B(n6121), .Z(n5467));
  OR2 U5955 ( .A(pi114), .B(n4885), .Z(n6120));
  AN2 U5956 ( .A(pi192), .B(n6122), .Z(n6113));
  OR2 U5957 ( .A(n6123), .B(n6124), .Z(n6122));
  AN2 U5958 ( .A(pi148), .B(n4881), .Z(n6124));
  AN2 U5959 ( .A(n4475), .B(n6125), .Z(n6123));
  OR2 U5960 ( .A(n5466), .B(n6126), .Z(n6125));
  IV2 U5961 ( .A(n5491), .Z(n6126));
  OR2 U5962 ( .A(po102), .B(n3901), .Z(n5491));
  IV2 U5963 ( .A(pi069), .Z(n3901));
  AN2 U5964 ( .A(n6127), .B(n6128), .Z(n5466));
  OR2 U5965 ( .A(pi069), .B(n4885), .Z(n6127));
  AN2 U5966 ( .A(n5461), .B(n4475), .Z(n6112));
  AN2 U5967 ( .A(n4087), .B(n6129), .Z(n5461));
  AN2 U5968 ( .A(n6130), .B(n4341), .Z(n6129));
  IV2 U5969 ( .A(n5474), .Z(n6130));
  AN2 U5970 ( .A(n6131), .B(po102), .Z(n5474));
  AN2 U5971 ( .A(n4334), .B(n4333), .Z(n4087));
  OR2 U5972 ( .A(n6132), .B(n4656), .Z(n4334));
  OR2 U5973 ( .A(n6133), .B(n6134), .Z(n4656));
  AN2 U5974 ( .A(n5074), .B(n3083), .Z(n6133));
  AN2 U5975 ( .A(n6135), .B(n3083), .Z(n6132));
  AN2 U5976 ( .A(n3018), .B(n4326), .Z(n6135));
  OR2 U5977 ( .A(n6136), .B(n5077), .Z(n4326));
  OR2 U5978 ( .A(n6137), .B(n3100), .Z(n5077));
  AN2 U5979 ( .A(n3280), .B(n4666), .Z(n6137));
  OR2 U5980 ( .A(n3286), .B(n6138), .Z(n4666));
  AN2 U5981 ( .A(n5829), .B(n3049), .Z(n3280));
  AN2 U5982 ( .A(n6139), .B(n3284), .Z(n6136));
  OR2 U5983 ( .A(n3049), .B(n5829), .Z(n3284));
  OR2 U5984 ( .A(n6140), .B(n3287), .Z(n6139));
  OR2 U5985 ( .A(n6141), .B(n6142), .Z(n3287));
  AN2 U5986 ( .A(pi141), .B(n3173), .Z(n6141));
  AN2 U5987 ( .A(n6143), .B(n3286), .Z(n6140));
  OR2 U5988 ( .A(n3173), .B(n3064), .Z(n6143));
  OR2 U5989 ( .A(n6144), .B(n6145), .Z(po000));
  AN2 U5990 ( .A(n6146), .B(po103), .Z(n6145));
  OR2 U5991 ( .A(n6147), .B(n6148), .Z(n6146));
  AN2 U5992 ( .A(n6149), .B(n3326), .Z(n6148));
  AN2 U5993 ( .A(n4217), .B(n3320), .Z(n6147));
  AN2 U5994 ( .A(n6150), .B(n3265), .Z(n6144));
  IV2 U5995 ( .A(po103), .Z(n3265));
  OR2 U5996 ( .A(n6151), .B(n6152), .Z(n6150));
  AN2 U5997 ( .A(n6149), .B(n3320), .Z(n6152));
  OR2 U5998 ( .A(n4406), .B(n4192), .Z(n3320));
  IV2 U5999 ( .A(n4205), .Z(n4192));
  AN2 U6000 ( .A(n4242), .B(n4331), .Z(n4406));
  IV2 U6001 ( .A(n4330), .Z(n4331));
  AN2 U6002 ( .A(n4217), .B(n3326), .Z(n6151));
  OR2 U6003 ( .A(n6153), .B(n4239), .Z(n3326));
  IV2 U6004 ( .A(n4242), .Z(n4239));
  OR2 U6005 ( .A(po028), .B(n6154), .Z(n4242));
  AN2 U6006 ( .A(n6155), .B(n6156), .Z(n6154));
  OR2 U6007 ( .A(n3321), .B(n3969), .Z(n6156));
  IV2 U6008 ( .A(pi169), .Z(n3969));
  AN2 U6009 ( .A(n4330), .B(n4205), .Z(n6153));
  OR2 U6010 ( .A(n6157), .B(n5056), .Z(n4205));
  IV2 U6011 ( .A(po028), .Z(n5056));
  AN2 U6012 ( .A(n3261), .B(n6158), .Z(n6157));
  OR2 U6013 ( .A(pi169), .B(n2837), .Z(n6158));
  OR2 U6014 ( .A(n6159), .B(n6160), .Z(n4330));
  OR2 U6015 ( .A(n6161), .B(n5930), .Z(n6160));
  OR2 U6016 ( .A(n6162), .B(n6163), .Z(n5930));
  OR2 U6017 ( .A(n6164), .B(n6165), .Z(n6163));
  AN2 U6018 ( .A(n3393), .B(n6166), .Z(n6165));
  OR2 U6019 ( .A(n6167), .B(n5853), .Z(n6166));
  AN2 U6020 ( .A(n6168), .B(n3371), .Z(n6167));
  IV2 U6021 ( .A(n3412), .Z(n3371));
  AN2 U6022 ( .A(n5999), .B(n6053), .Z(n6164));
  AN2 U6023 ( .A(n3453), .B(n3363), .Z(n5999));
  AN2 U6024 ( .A(n3926), .B(n4975), .Z(n6162));
  AN2 U6025 ( .A(n3940), .B(n4975), .Z(n6161));
  OR2 U6026 ( .A(n6169), .B(n6170), .Z(n6159));
  AN2 U6027 ( .A(n5931), .B(n6171), .Z(n6170));
  OR2 U6028 ( .A(n6172), .B(n6173), .Z(n6171));
  OR2 U6029 ( .A(n6174), .B(n6175), .Z(n6173));
  AN2 U6030 ( .A(n5888), .B(n3363), .Z(n6175));
  OR2 U6031 ( .A(n6176), .B(n6177), .Z(n5888));
  OR2 U6032 ( .A(n3248), .B(n6178), .Z(n6177));
  AN2 U6033 ( .A(n5833), .B(n3250), .Z(n6178));
  AN2 U6034 ( .A(n4937), .B(n6179), .Z(n5833));
  OR2 U6035 ( .A(n6180), .B(n6181), .Z(n6176));
  AN2 U6036 ( .A(n3495), .B(n5835), .Z(n6181));
  OR2 U6037 ( .A(n6182), .B(n5894), .Z(n5835));
  AN2 U6038 ( .A(n5966), .B(n6183), .Z(n6182));
  OR2 U6039 ( .A(n6184), .B(n6185), .Z(n5966));
  AN2 U6040 ( .A(pi171), .B(pi192), .Z(n6185));
  AN2 U6041 ( .A(pi142), .B(n2837), .Z(n6184));
  AN2 U6042 ( .A(n6186), .B(n5836), .Z(n6180));
  OR2 U6043 ( .A(n6187), .B(n6188), .Z(n5836));
  AN2 U6044 ( .A(n3705), .B(n5843), .Z(n6188));
  AN2 U6045 ( .A(pi192), .B(pi098), .Z(n3705));
  AN2 U6046 ( .A(n3717), .B(n6189), .Z(n6187));
  AN2 U6047 ( .A(n2837), .B(pi003), .Z(n3717));
  AN2 U6048 ( .A(n5889), .B(n3534), .Z(n6174));
  AN2 U6049 ( .A(n3261), .B(pi060), .Z(n3534));
  AN2 U6050 ( .A(pi192), .B(n6190), .Z(n5889));
  OR2 U6051 ( .A(n6191), .B(n6192), .Z(n6190));
  OR2 U6052 ( .A(n6193), .B(n6194), .Z(n6192));
  AN2 U6053 ( .A(pi004), .B(n4947), .Z(n6194));
  AN2 U6054 ( .A(n3640), .B(n3250), .Z(n6193));
  IV2 U6055 ( .A(n3344), .Z(n3250));
  IV2 U6056 ( .A(n3632), .Z(n3640));
  OR2 U6057 ( .A(po001), .B(n3998), .Z(n3632));
  OR2 U6058 ( .A(n6195), .B(n6196), .Z(n6191));
  AN2 U6059 ( .A(n6197), .B(n3495), .Z(n6196));
  AN2 U6060 ( .A(pi171), .B(n6183), .Z(n6197));
  AN2 U6061 ( .A(n6198), .B(n6186), .Z(n6195));
  IV2 U6062 ( .A(n6199), .Z(n6186));
  AN2 U6063 ( .A(pi098), .B(n5843), .Z(n6198));
  OR2 U6064 ( .A(pi171), .B(n4441), .Z(n5843));
  OR2 U6065 ( .A(n5892), .B(n6200), .Z(n6172));
  AN2 U6066 ( .A(n6201), .B(n5894), .Z(n6200));
  AN2 U6067 ( .A(n4441), .B(n4417), .Z(n5894));
  AN2 U6068 ( .A(n3495), .B(n3453), .Z(n6201));
  IV2 U6069 ( .A(n3451), .Z(n3453));
  OR2 U6070 ( .A(n3533), .B(n3321), .Z(n3451));
  IV2 U6071 ( .A(n3477), .Z(n3533));
  OR2 U6072 ( .A(pi060), .B(n2837), .Z(n3477));
  IV2 U6073 ( .A(n6202), .Z(n3495));
  IV2 U6074 ( .A(n6203), .Z(n5892));
  OR2 U6075 ( .A(n6204), .B(n6155), .Z(n6203));
  AN2 U6076 ( .A(n6205), .B(n6206), .Z(n6204));
  AN2 U6077 ( .A(n6207), .B(n6208), .Z(n6206));
  OR2 U6078 ( .A(n6199), .B(n6209), .Z(n6208));
  OR2 U6079 ( .A(n3244), .B(n3597), .Z(n6209));
  IV2 U6080 ( .A(pi003), .Z(n3597));
  IV2 U6081 ( .A(n6189), .Z(n3244));
  OR2 U6082 ( .A(pi142), .B(n4441), .Z(n6189));
  OR2 U6083 ( .A(n4418), .B(n6202), .Z(n6199));
  IV2 U6084 ( .A(n4426), .Z(n4418));
  OR2 U6085 ( .A(n3688), .B(n3290), .Z(n4426));
  IV2 U6086 ( .A(po011), .Z(n3688));
  OR2 U6087 ( .A(n6202), .B(n6210), .Z(n6207));
  OR2 U6088 ( .A(n4430), .B(n4440), .Z(n6210));
  IV2 U6089 ( .A(pi142), .Z(n4440));
  IV2 U6090 ( .A(n6183), .Z(n4430));
  OR2 U6091 ( .A(n4417), .B(n4441), .Z(n6183));
  IV2 U6092 ( .A(po036), .Z(n4441));
  IV2 U6093 ( .A(n3236), .Z(n4417));
  OR2 U6094 ( .A(n3234), .B(po011), .Z(n3236));
  IV2 U6095 ( .A(n3290), .Z(n3234));
  OR2 U6096 ( .A(n6211), .B(n6212), .Z(n3290));
  OR2 U6097 ( .A(n6213), .B(n6214), .Z(n6212));
  OR2 U6098 ( .A(n6215), .B(n6216), .Z(n6214));
  AN2 U6099 ( .A(pi192), .B(n5980), .Z(n6216));
  OR2 U6100 ( .A(n6217), .B(n6218), .Z(n5980));
  OR2 U6101 ( .A(n6219), .B(n6220), .Z(n6218));
  AN2 U6102 ( .A(pi045), .B(n4915), .Z(n6220));
  AN2 U6103 ( .A(n4621), .B(n4751), .Z(n6219));
  IV2 U6104 ( .A(n4465), .Z(n4621));
  OR2 U6105 ( .A(po014), .B(n3908), .Z(n4465));
  IV2 U6106 ( .A(pi079), .Z(n3908));
  OR2 U6107 ( .A(n6221), .B(n6222), .Z(n6217));
  AN2 U6108 ( .A(n6223), .B(n3757), .Z(n6222));
  AN2 U6109 ( .A(pi158), .B(n4628), .Z(n6223));
  AN2 U6110 ( .A(n6224), .B(n6225), .Z(n6221));
  AN2 U6111 ( .A(pi175), .B(n5037), .Z(n6224));
  AN2 U6112 ( .A(n6008), .B(n2837), .Z(n6215));
  OR2 U6113 ( .A(n6226), .B(n6227), .Z(n6008));
  OR2 U6114 ( .A(n6228), .B(n6229), .Z(n6227));
  AN2 U6115 ( .A(pi095), .B(n4915), .Z(n6229));
  AN2 U6116 ( .A(n4623), .B(n4751), .Z(n6228));
  IV2 U6117 ( .A(n4469), .Z(n4623));
  OR2 U6118 ( .A(po014), .B(n4648), .Z(n4469));
  IV2 U6119 ( .A(pi156), .Z(n4648));
  OR2 U6120 ( .A(n6230), .B(n6231), .Z(n6226));
  AN2 U6121 ( .A(n6232), .B(n3757), .Z(n6231));
  AN2 U6122 ( .A(pi151), .B(n4628), .Z(n6232));
  AN2 U6123 ( .A(n6233), .B(n6225), .Z(n6230));
  AN2 U6124 ( .A(pi185), .B(n5037), .Z(n6233));
  AN2 U6125 ( .A(n5985), .B(n6234), .Z(n6213));
  OR2 U6126 ( .A(n6235), .B(n6236), .Z(n6234));
  OR2 U6127 ( .A(n6237), .B(n6238), .Z(n6236));
  OR2 U6128 ( .A(n6239), .B(n6240), .Z(n6238));
  AN2 U6129 ( .A(n6241), .B(n3055), .Z(n6240));
  AN2 U6130 ( .A(n5822), .B(n3119), .Z(n6241));
  OR2 U6131 ( .A(n6242), .B(n6016), .Z(n3119));
  AN2 U6132 ( .A(pi141), .B(po099), .Z(n6242));
  AN2 U6133 ( .A(n5994), .B(n6243), .Z(n6239));
  AN2 U6134 ( .A(n6244), .B(n3049), .Z(n6237));
  OR2 U6135 ( .A(n6243), .B(n6245), .Z(n6244));
  OR2 U6136 ( .A(n6020), .B(n6246), .Z(n6245));
  AN2 U6137 ( .A(n6247), .B(n5826), .Z(n6246));
  AN2 U6138 ( .A(n3106), .B(n5829), .Z(n5826));
  OR2 U6139 ( .A(n5994), .B(n5822), .Z(n5829));
  IV2 U6140 ( .A(pi166), .Z(n3106));
  AN2 U6141 ( .A(n3063), .B(pi192), .Z(n6247));
  AN2 U6142 ( .A(n6016), .B(n5994), .Z(n6020));
  AN2 U6143 ( .A(n3286), .B(n3177), .Z(n6016));
  OR2 U6144 ( .A(n6142), .B(n6248), .Z(n6243));
  AN2 U6145 ( .A(n3207), .B(n3286), .Z(n6248));
  OR2 U6146 ( .A(n6249), .B(n6250), .Z(n3207));
  AN2 U6147 ( .A(n3064), .B(n3171), .Z(n6250));
  AN2 U6148 ( .A(n3173), .B(n3177), .Z(n6249));
  IV2 U6149 ( .A(pi141), .Z(n3177));
  AN2 U6150 ( .A(pi033), .B(n3064), .Z(n6142));
  OR2 U6151 ( .A(n6251), .B(n6252), .Z(n6235));
  OR2 U6152 ( .A(n6044), .B(n3100), .Z(n6252));
  AN2 U6153 ( .A(n3286), .B(n6138), .Z(n3100));
  OR2 U6154 ( .A(n6253), .B(n6254), .Z(n6138));
  AN2 U6155 ( .A(pi033), .B(pi192), .Z(n6254));
  AN2 U6156 ( .A(pi141), .B(n2837), .Z(n6253));
  AN2 U6157 ( .A(n6255), .B(pi141), .Z(n6044));
  OR2 U6158 ( .A(n3071), .B(n6256), .Z(n6255));
  AN2 U6159 ( .A(n3055), .B(n5994), .Z(n6256));
  IV2 U6160 ( .A(n6257), .Z(n5994));
  OR2 U6161 ( .A(n2925), .B(n5099), .Z(n6257));
  OR2 U6162 ( .A(n6258), .B(n6259), .Z(n5099));
  OR2 U6163 ( .A(n3146), .B(n6260), .Z(n6259));
  OR2 U6164 ( .A(n6261), .B(n6262), .Z(n6260));
  AN2 U6165 ( .A(n2845), .B(n2837), .Z(n6262));
  IV2 U6166 ( .A(n2846), .Z(n2845));
  AN2 U6167 ( .A(n6263), .B(n6264), .Z(n2846));
  OR2 U6168 ( .A(n3141), .B(po044), .Z(n6263));
  IV2 U6169 ( .A(pi201), .Z(n3141));
  AN2 U6170 ( .A(pi192), .B(n2833), .Z(n6261));
  IV2 U6171 ( .A(n2834), .Z(n2833));
  AN2 U6172 ( .A(n6265), .B(n6266), .Z(n2834));
  OR2 U6173 ( .A(n3136), .B(po044), .Z(n6265));
  IV2 U6174 ( .A(pi088), .Z(n3136));
  OR2 U6175 ( .A(n6267), .B(n6268), .Z(n3146));
  AN2 U6176 ( .A(n2880), .B(pi192), .Z(n6268));
  IV2 U6177 ( .A(n2878), .Z(n2880));
  OR2 U6178 ( .A(pi077), .B(n2962), .Z(n2878));
  AN2 U6179 ( .A(n2978), .B(n2837), .Z(n6267));
  IV2 U6180 ( .A(n2939), .Z(n2978));
  OR2 U6181 ( .A(n2998), .B(n6269), .Z(n6258));
  OR2 U6182 ( .A(n2901), .B(n2862), .Z(n6269));
  IV2 U6183 ( .A(pi200), .Z(n2901));
  IV2 U6184 ( .A(n3003), .Z(n2925));
  OR2 U6185 ( .A(pi192), .B(n2960), .Z(n3003));
  IV2 U6186 ( .A(n6270), .Z(n2960));
  OR2 U6187 ( .A(n6271), .B(n6272), .Z(n6270));
  AN2 U6188 ( .A(pi081), .B(n2931), .Z(n6272));
  IV2 U6189 ( .A(po107), .Z(n2931));
  AN2 U6190 ( .A(po107), .B(n2982), .Z(n6271));
  AN2 U6191 ( .A(n2837), .B(n6017), .Z(n3055));
  IV2 U6192 ( .A(n5828), .Z(n6017));
  OR2 U6193 ( .A(n6273), .B(n6015), .Z(n5828));
  AN2 U6194 ( .A(pi174), .B(n3049), .Z(n6015));
  AN2 U6195 ( .A(po010), .B(n5115), .Z(n6273));
  IV2 U6196 ( .A(pi174), .Z(n5115));
  AN2 U6197 ( .A(n3049), .B(n3173), .Z(n3071));
  AN2 U6198 ( .A(n2837), .B(pi174), .Z(n3173));
  IV2 U6199 ( .A(po010), .Z(n3049));
  AN2 U6200 ( .A(n6274), .B(n3063), .Z(n6251));
  IV2 U6201 ( .A(n6275), .Z(n3063));
  OR2 U6202 ( .A(n6276), .B(n6277), .Z(n6275));
  AN2 U6203 ( .A(pi033), .B(n3286), .Z(n6277));
  IV2 U6204 ( .A(po099), .Z(n3286));
  AN2 U6205 ( .A(po099), .B(n3171), .Z(n6276));
  IV2 U6206 ( .A(pi033), .Z(n3171));
  AN2 U6207 ( .A(n3064), .B(n5822), .Z(n6274));
  OR2 U6208 ( .A(n6278), .B(n6279), .Z(n5822));
  OR2 U6209 ( .A(n6280), .B(n6281), .Z(n6279));
  AN2 U6210 ( .A(n6282), .B(pi192), .Z(n6281));
  AN2 U6211 ( .A(n5156), .B(n6266), .Z(n6282));
  OR2 U6212 ( .A(pi088), .B(n5000), .Z(n6266));
  OR2 U6213 ( .A(n6283), .B(n5153), .Z(n5156));
  AN2 U6214 ( .A(n2861), .B(n6284), .Z(n6283));
  OR2 U6215 ( .A(n2885), .B(n2892), .Z(n6284));
  AN2 U6216 ( .A(n5008), .B(pi157), .Z(n2892));
  AN2 U6217 ( .A(n2930), .B(n2876), .Z(n2885));
  IV2 U6218 ( .A(n2887), .Z(n2876));
  OR2 U6219 ( .A(po031), .B(n3846), .Z(n2887));
  IV2 U6220 ( .A(pi077), .Z(n3846));
  AN2 U6221 ( .A(n6285), .B(n2837), .Z(n6280));
  AN2 U6222 ( .A(n5175), .B(n6264), .Z(n6285));
  OR2 U6223 ( .A(pi201), .B(n5000), .Z(n6264));
  OR2 U6224 ( .A(n6286), .B(n6287), .Z(n5175));
  AN2 U6225 ( .A(n2861), .B(n6288), .Z(n6286));
  OR2 U6226 ( .A(n6289), .B(n2929), .Z(n6288));
  IV2 U6227 ( .A(n2947), .Z(n2929));
  OR2 U6228 ( .A(po106), .B(n5431), .Z(n2947));
  IV2 U6229 ( .A(pi206), .Z(n5431));
  AN2 U6230 ( .A(n2930), .B(n4113), .Z(n6289));
  OR2 U6231 ( .A(n2919), .B(n2936), .Z(n4113));
  IV2 U6232 ( .A(n2946), .Z(n2936));
  OR2 U6233 ( .A(po031), .B(n2957), .Z(n2946));
  IV2 U6234 ( .A(pi082), .Z(n2957));
  AN2 U6235 ( .A(n2902), .B(n2939), .Z(n2919));
  OR2 U6236 ( .A(pi082), .B(n2962), .Z(n2939));
  IV2 U6237 ( .A(po031), .Z(n2962));
  IV2 U6238 ( .A(n2974), .Z(n2902));
  OR2 U6239 ( .A(po107), .B(n2982), .Z(n2974));
  IV2 U6240 ( .A(pi081), .Z(n2982));
  IV2 U6241 ( .A(n2862), .Z(n2930));
  OR2 U6242 ( .A(n6290), .B(n6291), .Z(n2862));
  AN2 U6243 ( .A(n6292), .B(n5008), .Z(n6291));
  IV2 U6244 ( .A(po106), .Z(n5008));
  AN2 U6245 ( .A(n6293), .B(po106), .Z(n6290));
  IV2 U6246 ( .A(n6292), .Z(n6293));
  OR2 U6247 ( .A(n6294), .B(n6295), .Z(n6292));
  AN2 U6248 ( .A(pi192), .B(pi157), .Z(n6295));
  AN2 U6249 ( .A(pi206), .B(n2837), .Z(n6294));
  IV2 U6250 ( .A(n2998), .Z(n2861));
  OR2 U6251 ( .A(n6296), .B(n6297), .Z(n2998));
  OR2 U6252 ( .A(n6298), .B(n6299), .Z(n6297));
  AN2 U6253 ( .A(n5153), .B(pi192), .Z(n6299));
  AN2 U6254 ( .A(n5004), .B(pi026), .Z(n5153));
  IV2 U6255 ( .A(po079), .Z(n5004));
  AN2 U6256 ( .A(n6287), .B(n2837), .Z(n6298));
  IV2 U6257 ( .A(n5172), .Z(n6287));
  OR2 U6258 ( .A(po079), .B(n5165), .Z(n5172));
  AN2 U6259 ( .A(po079), .B(n6027), .Z(n6296));
  OR2 U6260 ( .A(n6300), .B(n6301), .Z(n6027));
  AN2 U6261 ( .A(pi192), .B(n3847), .Z(n6301));
  IV2 U6262 ( .A(pi026), .Z(n3847));
  AN2 U6263 ( .A(n5165), .B(n2837), .Z(n6300));
  IV2 U6264 ( .A(pi107), .Z(n5165));
  AN2 U6265 ( .A(n3011), .B(n5000), .Z(n6278));
  IV2 U6266 ( .A(po044), .Z(n5000));
  OR2 U6267 ( .A(n6302), .B(n6303), .Z(n3011));
  AN2 U6268 ( .A(pi088), .B(pi192), .Z(n6303));
  AN2 U6269 ( .A(pi201), .B(n2837), .Z(n6302));
  AN2 U6270 ( .A(pi192), .B(pi166), .Z(n3064));
  AN2 U6271 ( .A(n3018), .B(n5984), .Z(n5985));
  AN2 U6272 ( .A(n6304), .B(n5104), .Z(n3018));
  IV2 U6273 ( .A(n5074), .Z(n5104));
  OR2 U6274 ( .A(n6305), .B(n5040), .Z(n6304));
  OR2 U6275 ( .A(n6306), .B(n6307), .Z(n6211));
  OR2 U6276 ( .A(n6308), .B(n6309), .Z(n6307));
  AN2 U6277 ( .A(n4624), .B(n5981), .Z(n6309));
  AN2 U6278 ( .A(n3300), .B(n3305), .Z(n4624));
  AN2 U6279 ( .A(n5984), .B(n5074), .Z(n6308));
  AN2 U6280 ( .A(n5040), .B(n6305), .Z(n5074));
  OR2 U6281 ( .A(n6310), .B(n6311), .Z(n6305));
  AN2 U6282 ( .A(pi096), .B(pi192), .Z(n6311));
  AN2 U6283 ( .A(pi128), .B(n2837), .Z(n6310));
  IV2 U6284 ( .A(po070), .Z(n5040));
  AN2 U6285 ( .A(n3083), .B(n6225), .Z(n5984));
  AN2 U6286 ( .A(n6312), .B(n6313), .Z(n6225));
  AN2 U6287 ( .A(n3760), .B(n4341), .Z(n6313));
  AN2 U6288 ( .A(n4333), .B(n4482), .Z(n6312));
  OR2 U6289 ( .A(n6314), .B(n6315), .Z(n4333));
  AN2 U6290 ( .A(po025), .B(n6316), .Z(n6315));
  OR2 U6291 ( .A(n6317), .B(n3888), .Z(n6316));
  AN2 U6292 ( .A(pi192), .B(pi191), .Z(n3888));
  AN2 U6293 ( .A(pi076), .B(n2837), .Z(n6317));
  AN2 U6294 ( .A(n3781), .B(n4557), .Z(n6314));
  OR2 U6295 ( .A(n4538), .B(n3890), .Z(n3781));
  IV2 U6296 ( .A(n6318), .Z(n3890));
  OR2 U6297 ( .A(pi191), .B(n2837), .Z(n6318));
  AN2 U6298 ( .A(n4077), .B(n2837), .Z(n4538));
  IV2 U6299 ( .A(n3021), .Z(n3083));
  OR2 U6300 ( .A(n6319), .B(n6134), .Z(n3021));
  AN2 U6301 ( .A(n6320), .B(n5037), .Z(n6134));
  IV2 U6302 ( .A(po035), .Z(n5037));
  AN2 U6303 ( .A(n6321), .B(po035), .Z(n6319));
  IV2 U6304 ( .A(n6320), .Z(n6321));
  OR2 U6305 ( .A(n6322), .B(n6323), .Z(n6320));
  AN2 U6306 ( .A(pi175), .B(pi192), .Z(n6323));
  AN2 U6307 ( .A(pi185), .B(n2837), .Z(n6322));
  AN2 U6308 ( .A(n3760), .B(n6324), .Z(n6306));
  OR2 U6309 ( .A(n6325), .B(n6326), .Z(n6324));
  OR2 U6310 ( .A(n6327), .B(n6328), .Z(n6326));
  AN2 U6311 ( .A(n4482), .B(n4340), .Z(n6328));
  OR2 U6312 ( .A(n6329), .B(n6330), .Z(n4340));
  AN2 U6313 ( .A(n6121), .B(n2837), .Z(n6330));
  OR2 U6314 ( .A(n6331), .B(n4567), .Z(n6121));
  IV2 U6315 ( .A(n4578), .Z(n4567));
  OR2 U6316 ( .A(po024), .B(n4358), .Z(n4578));
  AN2 U6317 ( .A(n4084), .B(n4066), .Z(n6331));
  OR2 U6318 ( .A(n6332), .B(n4539), .Z(n4084));
  IV2 U6319 ( .A(n5503), .Z(n4539));
  OR2 U6320 ( .A(po059), .B(n4074), .Z(n5503));
  IV2 U6321 ( .A(pi170), .Z(n4074));
  AN2 U6322 ( .A(n4576), .B(n3778), .Z(n6332));
  IV2 U6323 ( .A(n4580), .Z(n4576));
  OR2 U6324 ( .A(po025), .B(n4077), .Z(n4580));
  IV2 U6325 ( .A(pi076), .Z(n4077));
  AN2 U6326 ( .A(pi192), .B(n6128), .Z(n6329));
  OR2 U6327 ( .A(n6333), .B(n6334), .Z(n6128));
  OR2 U6328 ( .A(n4561), .B(n6335), .Z(n6334));
  AN2 U6329 ( .A(n6336), .B(n4341), .Z(n6335));
  AN2 U6330 ( .A(n4066), .B(n3778), .Z(n4341));
  IV2 U6331 ( .A(n3773), .Z(n3778));
  OR2 U6332 ( .A(n6337), .B(n6338), .Z(n3773));
  AN2 U6333 ( .A(n6339), .B(n4877), .Z(n6338));
  IV2 U6334 ( .A(po059), .Z(n4877));
  AN2 U6335 ( .A(n6340), .B(po059), .Z(n6337));
  IV2 U6336 ( .A(n6339), .Z(n6340));
  OR2 U6337 ( .A(n6341), .B(n6342), .Z(n6339));
  AN2 U6338 ( .A(pi135), .B(pi192), .Z(n6342));
  AN2 U6339 ( .A(pi170), .B(n2837), .Z(n6341));
  AN2 U6340 ( .A(pi191), .B(n4557), .Z(n6336));
  IV2 U6341 ( .A(po025), .Z(n4557));
  IV2 U6342 ( .A(n4348), .Z(n4561));
  OR2 U6343 ( .A(po024), .B(n3896), .Z(n4348));
  AN2 U6344 ( .A(n4085), .B(n4066), .Z(n6333));
  OR2 U6345 ( .A(n6343), .B(n6344), .Z(n4066));
  OR2 U6346 ( .A(n6345), .B(n6346), .Z(n6344));
  AN2 U6347 ( .A(n6347), .B(po024), .Z(n6346));
  AN2 U6348 ( .A(pi005), .B(pi192), .Z(n6347));
  AN2 U6349 ( .A(n6348), .B(n4874), .Z(n6345));
  IV2 U6350 ( .A(po024), .Z(n4874));
  OR2 U6351 ( .A(n6349), .B(n5483), .Z(n6348));
  AN2 U6352 ( .A(pi192), .B(n3896), .Z(n5483));
  IV2 U6353 ( .A(pi005), .Z(n3896));
  AN2 U6354 ( .A(n4358), .B(n2837), .Z(n6349));
  IV2 U6355 ( .A(pi160), .Z(n4358));
  AN2 U6356 ( .A(pi160), .B(n5477), .Z(n6343));
  AN2 U6357 ( .A(n2837), .B(po024), .Z(n5477));
  IV2 U6358 ( .A(n4353), .Z(n4085));
  OR2 U6359 ( .A(po059), .B(n3880), .Z(n4353));
  IV2 U6360 ( .A(pi135), .Z(n3880));
  AN2 U6361 ( .A(n4342), .B(n4475), .Z(n4482));
  AN2 U6362 ( .A(n6350), .B(n6351), .Z(n4342));
  OR2 U6363 ( .A(n6131), .B(po102), .Z(n6351));
  IV2 U6364 ( .A(n6352), .Z(n6131));
  OR2 U6365 ( .A(n6352), .B(n4885), .Z(n6350));
  AN2 U6366 ( .A(n5462), .B(n4475), .Z(n6327));
  IV2 U6367 ( .A(n4478), .Z(n4475));
  OR2 U6368 ( .A(n6353), .B(n6325), .Z(n4478));
  AN2 U6369 ( .A(n6354), .B(po072), .Z(n6353));
  IV2 U6370 ( .A(n6355), .Z(n6354));
  AN2 U6371 ( .A(n6352), .B(n4885), .Z(n5462));
  IV2 U6372 ( .A(po102), .Z(n4885));
  OR2 U6373 ( .A(n6356), .B(n6357), .Z(n6352));
  AN2 U6374 ( .A(pi069), .B(pi192), .Z(n6357));
  AN2 U6375 ( .A(pi114), .B(n2837), .Z(n6356));
  AN2 U6376 ( .A(n6355), .B(n4881), .Z(n6325));
  IV2 U6377 ( .A(po072), .Z(n4881));
  OR2 U6378 ( .A(n6358), .B(n6359), .Z(n6355));
  AN2 U6379 ( .A(pi148), .B(pi192), .Z(n6359));
  AN2 U6380 ( .A(pi108), .B(n2837), .Z(n6358));
  AN2 U6381 ( .A(n4450), .B(n5981), .Z(n3760));
  AN2 U6382 ( .A(n3301), .B(n4751), .Z(n5981));
  AN2 U6383 ( .A(n4006), .B(n3757), .Z(n4751));
  IV2 U6384 ( .A(n4444), .Z(n3757));
  OR2 U6385 ( .A(n6360), .B(n3754), .Z(n4444));
  AN2 U6386 ( .A(n6361), .B(n4915), .Z(n3754));
  IV2 U6387 ( .A(po063), .Z(n4915));
  AN2 U6388 ( .A(n6362), .B(po063), .Z(n6360));
  IV2 U6389 ( .A(n6361), .Z(n6362));
  OR2 U6390 ( .A(n6363), .B(n6364), .Z(n6361));
  AN2 U6391 ( .A(pi045), .B(pi192), .Z(n6364));
  AN2 U6392 ( .A(pi095), .B(n2837), .Z(n6363));
  AN2 U6393 ( .A(n6365), .B(n6366), .Z(n4006));
  OR2 U6394 ( .A(n6367), .B(po092), .Z(n6366));
  IV2 U6395 ( .A(n4752), .Z(n6367));
  OR2 U6396 ( .A(n4752), .B(n4628), .Z(n6365));
  IV2 U6397 ( .A(po092), .Z(n4628));
  OR2 U6398 ( .A(n6368), .B(n6369), .Z(n4752));
  AN2 U6399 ( .A(pi158), .B(pi192), .Z(n6369));
  AN2 U6400 ( .A(pi151), .B(n2837), .Z(n6368));
  IV2 U6401 ( .A(n3295), .Z(n3301));
  OR2 U6402 ( .A(n6370), .B(n6371), .Z(n3295));
  AN2 U6403 ( .A(n4703), .B(n4861), .Z(n6371));
  IV2 U6404 ( .A(po014), .Z(n4861));
  AN2 U6405 ( .A(n4736), .B(po014), .Z(n6370));
  IV2 U6406 ( .A(n4703), .Z(n4736));
  OR2 U6407 ( .A(n6372), .B(n6373), .Z(n4703));
  AN2 U6408 ( .A(pi079), .B(pi192), .Z(n6373));
  AN2 U6409 ( .A(pi156), .B(n2837), .Z(n6372));
  IV2 U6410 ( .A(n4606), .Z(n4450));
  AN2 U6411 ( .A(n6374), .B(n6375), .Z(n4606));
  OR2 U6412 ( .A(n3305), .B(po039), .Z(n6375));
  OR2 U6413 ( .A(n3300), .B(n6376), .Z(n6374));
  IV2 U6414 ( .A(n3305), .Z(n6376));
  OR2 U6415 ( .A(n4685), .B(n4692), .Z(n3305));
  AN2 U6416 ( .A(pi192), .B(pi016), .Z(n4692));
  AN2 U6417 ( .A(n2837), .B(pi040), .Z(n4685));
  IV2 U6418 ( .A(po039), .Z(n3300));
  OR2 U6419 ( .A(n3352), .B(n3344), .Z(n6202));
  AN2 U6420 ( .A(n6377), .B(n6378), .Z(n3352));
  OR2 U6421 ( .A(n6179), .B(po001), .Z(n6378));
  IV2 U6422 ( .A(n6379), .Z(n6179));
  OR2 U6423 ( .A(n6379), .B(n4937), .Z(n6377));
  IV2 U6424 ( .A(po001), .Z(n4937));
  OR2 U6425 ( .A(n5959), .B(n6380), .Z(n6379));
  AN2 U6426 ( .A(pi192), .B(n3998), .Z(n6380));
  IV2 U6427 ( .A(pi068), .Z(n3998));
  AN2 U6428 ( .A(n2837), .B(n5379), .Z(n5959));
  AN2 U6429 ( .A(n6381), .B(n6382), .Z(n6205));
  OR2 U6430 ( .A(n3344), .B(n3590), .Z(n6382));
  OR2 U6431 ( .A(po001), .B(n5379), .Z(n3590));
  IV2 U6432 ( .A(pi195), .Z(n5379));
  OR2 U6433 ( .A(n6383), .B(n3248), .Z(n3344));
  AN2 U6434 ( .A(n6384), .B(n4947), .Z(n3248));
  IV2 U6435 ( .A(po082), .Z(n4947));
  AN2 U6436 ( .A(n6385), .B(po082), .Z(n6383));
  IV2 U6437 ( .A(n6384), .Z(n6385));
  OR2 U6438 ( .A(n6386), .B(n6387), .Z(n6384));
  AN2 U6439 ( .A(pi004), .B(pi192), .Z(n6387));
  AN2 U6440 ( .A(pi130), .B(n2837), .Z(n6386));
  OR2 U6441 ( .A(po082), .B(n5372), .Z(n6381));
  IV2 U6442 ( .A(pi130), .Z(n5372));
  AN2 U6443 ( .A(n3225), .B(n6053), .Z(n5931));
  IV2 U6444 ( .A(n3247), .Z(n3225));
  OR2 U6445 ( .A(n6388), .B(n3490), .Z(n3247));
  AN2 U6446 ( .A(n4943), .B(n5895), .Z(n3490));
  OR2 U6447 ( .A(n3926), .B(n3989), .Z(n5895));
  IV2 U6448 ( .A(n6389), .Z(n6388));
  OR2 U6449 ( .A(n4943), .B(n6390), .Z(n6389));
  AN2 U6450 ( .A(n6391), .B(n3261), .Z(n6390));
  OR2 U6451 ( .A(n2837), .B(pi133), .Z(n6391));
  AN2 U6452 ( .A(n6392), .B(n6053), .Z(n6169));
  AN2 U6453 ( .A(n3393), .B(n6393), .Z(n6053));
  IV2 U6454 ( .A(n3461), .Z(n6393));
  OR2 U6455 ( .A(n3401), .B(n3412), .Z(n3461));
  OR2 U6456 ( .A(n6394), .B(n5853), .Z(n3412));
  OR2 U6457 ( .A(n3466), .B(n3392), .Z(n5853));
  AN2 U6458 ( .A(n3380), .B(n3926), .Z(n3392));
  IV2 U6459 ( .A(po071), .Z(n3380));
  AN2 U6460 ( .A(n3261), .B(n3381), .Z(n3466));
  IV2 U6461 ( .A(n3399), .Z(n3381));
  OR2 U6462 ( .A(po071), .B(n3913), .Z(n3399));
  AN2 U6463 ( .A(po071), .B(n5878), .Z(n6394));
  OR2 U6464 ( .A(n3480), .B(n3321), .Z(n5878));
  AN2 U6465 ( .A(n3913), .B(pi192), .Z(n3480));
  IV2 U6466 ( .A(pi118), .Z(n3913));
  OR2 U6467 ( .A(n5881), .B(n6395), .Z(n3401));
  OR2 U6468 ( .A(n6168), .B(n6396), .Z(n6395));
  AN2 U6469 ( .A(po104), .B(n3321), .Z(n6396));
  AN2 U6470 ( .A(n3485), .B(n3261), .Z(n6168));
  IV2 U6471 ( .A(n3419), .Z(n3485));
  OR2 U6472 ( .A(n6397), .B(po104), .Z(n3419));
  AN2 U6473 ( .A(pi192), .B(n3942), .Z(n6397));
  IV2 U6474 ( .A(pi196), .Z(n3942));
  AN2 U6475 ( .A(pi192), .B(n5872), .Z(n5881));
  IV2 U6476 ( .A(n5866), .Z(n5872));
  OR2 U6477 ( .A(pi196), .B(n3512), .Z(n5866));
  IV2 U6478 ( .A(po104), .Z(n3512));
  OR2 U6479 ( .A(n6398), .B(n6399), .Z(n3393));
  AN2 U6480 ( .A(n6400), .B(n4975), .Z(n6399));
  IV2 U6481 ( .A(po038), .Z(n4975));
  OR2 U6482 ( .A(n6401), .B(n3321), .Z(n6400));
  AN2 U6483 ( .A(pi192), .B(n3943), .Z(n6401));
  IV2 U6484 ( .A(pi050), .Z(n3943));
  AN2 U6485 ( .A(po038), .B(n6402), .Z(n6398));
  OR2 U6486 ( .A(n3940), .B(n3926), .Z(n6402));
  AN2 U6487 ( .A(n3261), .B(pi050), .Z(n3940));
  AN2 U6488 ( .A(n6403), .B(n4943), .Z(n6392));
  IV2 U6489 ( .A(po057), .Z(n4943));
  OR2 U6490 ( .A(n6404), .B(n6052), .Z(n6403));
  OR2 U6491 ( .A(n6405), .B(n3926), .Z(n6052));
  IV2 U6492 ( .A(n6155), .Z(n3926));
  OR2 U6493 ( .A(pi192), .B(n3321), .Z(n6155));
  AN2 U6494 ( .A(pi060), .B(n3989), .Z(n6405));
  AN2 U6495 ( .A(n3989), .B(n3363), .Z(n6404));
  IV2 U6496 ( .A(po027), .Z(n3363));
  AN2 U6497 ( .A(n3261), .B(pi133), .Z(n3989));
  IV2 U6498 ( .A(n3321), .Z(n3261));
  IV2 U6499 ( .A(n6149), .Z(n4217));
  OR2 U6500 ( .A(n4148), .B(n3321), .Z(n6149));
  AN2 U6501 ( .A(pi161), .B(pi012), .Z(n3321));
  IV2 U6502 ( .A(n4247), .Z(n4148));
  OR2 U6503 ( .A(pi058), .B(n2837), .Z(n4247));
  IV2 U6504 ( .A(pi192), .Z(n2837));

endmodule

module IV2(A,  Z);
  input A;
  output Z;

  assign Z = ~A;
endmodule

module AN2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A & B;
endmodule

module OR2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A | B;
endmodule
