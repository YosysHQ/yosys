module test(input in, output out);
//no buffer removal
assign out = in;
endmodule
