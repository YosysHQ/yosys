// ---------------------------------------

module \$__ABC9_DPR16X4_COMB (input [3:0] $DO, RAD, output [3:0] DO);
    assign DO = $DO;
endmodule
