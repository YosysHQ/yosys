module test (y);
    output signed [2:0] y = 1'bf;
endmodule
