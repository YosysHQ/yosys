module \$__MISTRAL_MLAB (PORT_W_CLK, PORT_W_ADDR, PORT_W_WR_DATA, PORT_W_WR_EN, PORT_R_ADDR, PORT_R_RD_DATA);

parameter INIT = 0;

input PORT_W_CLK;
input [4:0] PORT_W_ADDR, PORT_R_ADDR;
input [4:0] PORT_W_WR_DATA;
input PORT_W_WR_EN;
output reg PORT_R_RD_DATA;

MISTRAL_MLAB _TECHMAP_REPLACE_ (.CLK1(PORT_W_CLK), .A1ADDR(PORT_W_ADDR), .A1DATA(PORT_W_WR_DATA), .A1EN(PORT_W_WR_EN), .B1ADDR(PORT_R_ADDR), .B1DATA(PORT_R_RD_DATA));

endmodule
