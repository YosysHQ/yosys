`ifdef INIT_LOWER
.INIT_00(permute_init(INIT[  0*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_01(permute_init(INIT[  1*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_02(permute_init(INIT[  2*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_03(permute_init(INIT[  3*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_04(permute_init(INIT[  4*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_05(permute_init(INIT[  5*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_06(permute_init(INIT[  6*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_07(permute_init(INIT[  7*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_08(permute_init(INIT[  8*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_09(permute_init(INIT[  9*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0A(permute_init(INIT[ 10*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0B(permute_init(INIT[ 11*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0C(permute_init(INIT[ 12*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0D(permute_init(INIT[ 13*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0E(permute_init(INIT[ 14*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0F(permute_init(INIT[ 15*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_10(permute_init(INIT[ 16*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_11(permute_init(INIT[ 17*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_12(permute_init(INIT[ 18*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_13(permute_init(INIT[ 19*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_14(permute_init(INIT[ 20*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_15(permute_init(INIT[ 21*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_16(permute_init(INIT[ 22*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_17(permute_init(INIT[ 23*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_18(permute_init(INIT[ 24*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_19(permute_init(INIT[ 25*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1A(permute_init(INIT[ 26*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1B(permute_init(INIT[ 27*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1C(permute_init(INIT[ 28*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1D(permute_init(INIT[ 29*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1E(permute_init(INIT[ 30*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1F(permute_init(INIT[ 31*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_20(permute_init(INIT[ 32*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_21(permute_init(INIT[ 33*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_22(permute_init(INIT[ 34*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_23(permute_init(INIT[ 35*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_24(permute_init(INIT[ 36*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_25(permute_init(INIT[ 37*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_26(permute_init(INIT[ 38*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_27(permute_init(INIT[ 39*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_28(permute_init(INIT[ 40*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_29(permute_init(INIT[ 41*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2A(permute_init(INIT[ 42*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2B(permute_init(INIT[ 43*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2C(permute_init(INIT[ 44*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2D(permute_init(INIT[ 45*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2E(permute_init(INIT[ 46*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2F(permute_init(INIT[ 47*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_30(permute_init(INIT[ 48*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_31(permute_init(INIT[ 49*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_32(permute_init(INIT[ 50*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_33(permute_init(INIT[ 51*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_34(permute_init(INIT[ 52*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_35(permute_init(INIT[ 53*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_36(permute_init(INIT[ 54*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_37(permute_init(INIT[ 55*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_38(permute_init(INIT[ 56*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_39(permute_init(INIT[ 57*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3A(permute_init(INIT[ 58*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3B(permute_init(INIT[ 59*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3C(permute_init(INIT[ 60*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3D(permute_init(INIT[ 61*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3E(permute_init(INIT[ 62*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3F(permute_init(INIT[ 63*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_40(permute_init(INIT[ 64*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_41(permute_init(INIT[ 65*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_42(permute_init(INIT[ 66*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_43(permute_init(INIT[ 67*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_44(permute_init(INIT[ 68*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_45(permute_init(INIT[ 69*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_46(permute_init(INIT[ 70*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_47(permute_init(INIT[ 71*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_48(permute_init(INIT[ 72*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_49(permute_init(INIT[ 73*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4A(permute_init(INIT[ 74*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4B(permute_init(INIT[ 75*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4C(permute_init(INIT[ 76*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4D(permute_init(INIT[ 77*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4E(permute_init(INIT[ 78*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4F(permute_init(INIT[ 79*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_50(permute_init(INIT[ 80*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_51(permute_init(INIT[ 81*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_52(permute_init(INIT[ 82*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_53(permute_init(INIT[ 83*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_54(permute_init(INIT[ 84*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_55(permute_init(INIT[ 85*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_56(permute_init(INIT[ 86*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_57(permute_init(INIT[ 87*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_58(permute_init(INIT[ 88*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_59(permute_init(INIT[ 89*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5A(permute_init(INIT[ 90*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5B(permute_init(INIT[ 91*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5C(permute_init(INIT[ 92*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5D(permute_init(INIT[ 93*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5E(permute_init(INIT[ 94*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5F(permute_init(INIT[ 95*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_60(permute_init(INIT[ 96*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_61(permute_init(INIT[ 97*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_62(permute_init(INIT[ 98*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_63(permute_init(INIT[ 99*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_64(permute_init(INIT[100*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_65(permute_init(INIT[101*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_66(permute_init(INIT[102*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_67(permute_init(INIT[103*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_68(permute_init(INIT[104*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_69(permute_init(INIT[105*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6A(permute_init(INIT[106*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6B(permute_init(INIT[107*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6C(permute_init(INIT[108*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6D(permute_init(INIT[109*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6E(permute_init(INIT[110*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6F(permute_init(INIT[111*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_70(permute_init(INIT[112*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_71(permute_init(INIT[113*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_72(permute_init(INIT[114*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_73(permute_init(INIT[115*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_74(permute_init(INIT[116*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_75(permute_init(INIT[117*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_76(permute_init(INIT[118*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_77(permute_init(INIT[119*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_78(permute_init(INIT[120*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_79(permute_init(INIT[121*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7A(permute_init(INIT[122*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7B(permute_init(INIT[123*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7C(permute_init(INIT[124*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7D(permute_init(INIT[125*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7E(permute_init(INIT[126*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7F(permute_init(INIT[127*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
`endif
`ifdef INIT_UPPER
.INIT_00(permute_init(INIT[128*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_01(permute_init(INIT[129*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_02(permute_init(INIT[130*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_03(permute_init(INIT[131*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_04(permute_init(INIT[132*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_05(permute_init(INIT[133*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_06(permute_init(INIT[134*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_07(permute_init(INIT[135*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_08(permute_init(INIT[136*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_09(permute_init(INIT[137*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0A(permute_init(INIT[138*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0B(permute_init(INIT[139*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0C(permute_init(INIT[140*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0D(permute_init(INIT[141*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0E(permute_init(INIT[142*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_0F(permute_init(INIT[143*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_10(permute_init(INIT[144*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_11(permute_init(INIT[145*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_12(permute_init(INIT[146*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_13(permute_init(INIT[147*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_14(permute_init(INIT[148*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_15(permute_init(INIT[149*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_16(permute_init(INIT[150*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_17(permute_init(INIT[151*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_18(permute_init(INIT[152*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_19(permute_init(INIT[153*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1A(permute_init(INIT[154*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1B(permute_init(INIT[155*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1C(permute_init(INIT[156*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1D(permute_init(INIT[157*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1E(permute_init(INIT[158*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_1F(permute_init(INIT[159*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_20(permute_init(INIT[160*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_21(permute_init(INIT[161*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_22(permute_init(INIT[162*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_23(permute_init(INIT[163*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_24(permute_init(INIT[164*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_25(permute_init(INIT[165*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_26(permute_init(INIT[166*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_27(permute_init(INIT[167*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_28(permute_init(INIT[168*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_29(permute_init(INIT[169*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2A(permute_init(INIT[170*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2B(permute_init(INIT[171*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2C(permute_init(INIT[172*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2D(permute_init(INIT[173*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2E(permute_init(INIT[174*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_2F(permute_init(INIT[175*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_30(permute_init(INIT[176*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_31(permute_init(INIT[177*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_32(permute_init(INIT[178*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_33(permute_init(INIT[179*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_34(permute_init(INIT[180*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_35(permute_init(INIT[181*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_36(permute_init(INIT[182*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_37(permute_init(INIT[183*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_38(permute_init(INIT[184*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_39(permute_init(INIT[185*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3A(permute_init(INIT[186*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3B(permute_init(INIT[187*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3C(permute_init(INIT[188*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3D(permute_init(INIT[189*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3E(permute_init(INIT[190*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_3F(permute_init(INIT[191*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_40(permute_init(INIT[192*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_41(permute_init(INIT[193*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_42(permute_init(INIT[194*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_43(permute_init(INIT[195*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_44(permute_init(INIT[196*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_45(permute_init(INIT[197*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_46(permute_init(INIT[198*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_47(permute_init(INIT[199*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_48(permute_init(INIT[200*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_49(permute_init(INIT[201*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4A(permute_init(INIT[202*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4B(permute_init(INIT[203*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4C(permute_init(INIT[204*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4D(permute_init(INIT[205*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4E(permute_init(INIT[206*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_4F(permute_init(INIT[207*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_50(permute_init(INIT[208*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_51(permute_init(INIT[209*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_52(permute_init(INIT[210*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_53(permute_init(INIT[211*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_54(permute_init(INIT[212*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_55(permute_init(INIT[213*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_56(permute_init(INIT[214*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_57(permute_init(INIT[215*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_58(permute_init(INIT[216*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_59(permute_init(INIT[217*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5A(permute_init(INIT[218*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5B(permute_init(INIT[219*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5C(permute_init(INIT[220*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5D(permute_init(INIT[221*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5E(permute_init(INIT[222*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_5F(permute_init(INIT[223*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_60(permute_init(INIT[224*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_61(permute_init(INIT[225*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_62(permute_init(INIT[226*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_63(permute_init(INIT[227*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_64(permute_init(INIT[228*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_65(permute_init(INIT[229*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_66(permute_init(INIT[230*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_67(permute_init(INIT[231*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_68(permute_init(INIT[232*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_69(permute_init(INIT[233*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6A(permute_init(INIT[234*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6B(permute_init(INIT[235*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6C(permute_init(INIT[236*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6D(permute_init(INIT[237*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6E(permute_init(INIT[238*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_6F(permute_init(INIT[239*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_70(permute_init(INIT[240*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_71(permute_init(INIT[241*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_72(permute_init(INIT[242*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_73(permute_init(INIT[243*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_74(permute_init(INIT[244*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_75(permute_init(INIT[245*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_76(permute_init(INIT[246*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_77(permute_init(INIT[247*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_78(permute_init(INIT[248*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_79(permute_init(INIT[249*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7A(permute_init(INIT[250*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7B(permute_init(INIT[251*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7C(permute_init(INIT[252*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7D(permute_init(INIT[253*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7E(permute_init(INIT[254*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
.INIT_7F(permute_init(INIT[255*INIT_CHUNK_SIZE +: INIT_CHUNK_SIZE])),
`endif
