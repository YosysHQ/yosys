module typedef_test;
  typedef integer intA;
  typedef reg [31:0] word;
  typedef word fourbytes;
  intA a;
  word w;
  fourbytes f;
endmodule
