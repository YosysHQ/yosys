module test(input in, output  out);

assign out = -in;

endmodule
