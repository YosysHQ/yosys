module a;
initial
begin : label1
end: label2
endmodule

