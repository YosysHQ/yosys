module my_module(
		 input	a,
		 input	b,
		 output	sum
		 );
   // Perform addition
   assign sum = a + b;

endmodule
