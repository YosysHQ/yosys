(* blackbox *)
module ACC84_2DSP(clk, rst, X, Z);
    input [83:0] X;
    output [84:0] Z;
    input clk;
    input rst;
    parameter g_pipe = 2;
endmodule

(* blackbox *)
module ACC92_2DSP(clk, rst, X, Z);
    input [55:0] X;
    output [91:0] Z;
    input clk;
    input rst;
    parameter g_pipe = 2;
endmodule

(* blackbox *)
module ACC98_2DSP(clk, rst, X, Z);
    input [55:0] X;
    output [97:0] Z;
    input clk;
    input rst;
    parameter g_pipe = 2;
endmodule

(* blackbox *)
module ADD84_1DSP_2CYCLES(clk, rst, X, Y, Z);
    input [41:0] X;
    input [41:0] Y;
    output [84:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module ADD84_2DSP(clk, rst, X, Y, Z);
    input [83:0] X;
    input [83:0] Y;
    output [84:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module NX_BD(I, O);
    input I;
    output O;
    parameter mode = "global_lowskew";
endmodule

(* blackbox *)
module NX_BFF(I, O);
    input I;
    output O;
endmodule

(* blackbox *)
module NX_BFR(I, O);
    input I;
    output O;
    parameter data_inv = 1'b0;
    parameter iobname = "";
    parameter location = "";
    parameter mode = 0;
    parameter path = 0;
    parameter ring = 0;
endmodule

(* blackbox *)
module NX_CRX_L(DSCR_E_I, DEC_E_I, ALIGN_E_I, ALIGN_S_I, REP_E_I, BUF_R_I, OVS_BS_I1, OVS_BS_I2, BUF_FE_I, RST_N_I, CDR_R_I, CKG_RN_I, PLL_RN_I, TST_I1, TST_I2, TST_I3, TST_I4, LOS_O, DATA_O1, DATA_O2, DATA_O3
, DATA_O4, DATA_O5, DATA_O6, DATA_O7, DATA_O8, DATA_O9, DATA_O10, DATA_O11, DATA_O12, DATA_O13, DATA_O14, DATA_O15, DATA_O16, DATA_O17, DATA_O18, DATA_O19, DATA_O20, DATA_O21, DATA_O22, DATA_O23, DATA_O24
, DATA_O25, DATA_O26, DATA_O27, DATA_O28, DATA_O29, DATA_O30, DATA_O31, DATA_O32, DATA_O33, DATA_O34, DATA_O35, DATA_O36, DATA_O37, DATA_O38, DATA_O39, DATA_O40, DATA_O41, DATA_O42, DATA_O43, DATA_O44, DATA_O45
, DATA_O46, DATA_O47, DATA_O48, DATA_O49, DATA_O50, DATA_O51, DATA_O52, DATA_O53, DATA_O54, DATA_O55, DATA_O56, DATA_O57, DATA_O58, DATA_O59, DATA_O60, DATA_O61, DATA_O62, DATA_O63, DATA_O64, CH_COM_O1, CH_COM_O2
, CH_COM_O3, CH_COM_O4, CH_COM_O5, CH_COM_O6, CH_COM_O7, CH_COM_O8, CH_K_O1, CH_K_O2, CH_K_O3, CH_K_O4, CH_K_O5, CH_K_O6, CH_K_O7, CH_K_O8, NIT_O1, NIT_O2, NIT_O3, NIT_O4, NIT_O5, NIT_O6, NIT_O7
, NIT_O8, D_ERR_O1, D_ERR_O2, D_ERR_O3, D_ERR_O4, D_ERR_O5, D_ERR_O6, D_ERR_O7, D_ERR_O8, CH_A_O1, CH_A_O2, CH_A_O3, CH_A_O4, CH_A_O5, CH_A_O6, CH_A_O7, CH_A_O8, CH_F_O1, CH_F_O2, CH_F_O3, CH_F_O4
, CH_F_O5, CH_F_O6, CH_F_O7, CH_F_O8, ALIGN_O, BUSY_O, TST_O1, TST_O2, TST_O3, TST_O4, TST_O5, TST_O6, TST_O7, TST_O8, LOCK_O, RX_I, LINK);
    input ALIGN_E_I;
    output ALIGN_O;
    input ALIGN_S_I;
    input BUF_FE_I;
    input BUF_R_I;
    output BUSY_O;
    input CDR_R_I;
    output CH_A_O1;
    output CH_A_O2;
    output CH_A_O3;
    output CH_A_O4;
    output CH_A_O5;
    output CH_A_O6;
    output CH_A_O7;
    output CH_A_O8;
    output CH_COM_O1;
    output CH_COM_O2;
    output CH_COM_O3;
    output CH_COM_O4;
    output CH_COM_O5;
    output CH_COM_O6;
    output CH_COM_O7;
    output CH_COM_O8;
    output CH_F_O1;
    output CH_F_O2;
    output CH_F_O3;
    output CH_F_O4;
    output CH_F_O5;
    output CH_F_O6;
    output CH_F_O7;
    output CH_F_O8;
    output CH_K_O1;
    output CH_K_O2;
    output CH_K_O3;
    output CH_K_O4;
    output CH_K_O5;
    output CH_K_O6;
    output CH_K_O7;
    output CH_K_O8;
    input CKG_RN_I;
    output DATA_O1;
    output DATA_O10;
    output DATA_O11;
    output DATA_O12;
    output DATA_O13;
    output DATA_O14;
    output DATA_O15;
    output DATA_O16;
    output DATA_O17;
    output DATA_O18;
    output DATA_O19;
    output DATA_O2;
    output DATA_O20;
    output DATA_O21;
    output DATA_O22;
    output DATA_O23;
    output DATA_O24;
    output DATA_O25;
    output DATA_O26;
    output DATA_O27;
    output DATA_O28;
    output DATA_O29;
    output DATA_O3;
    output DATA_O30;
    output DATA_O31;
    output DATA_O32;
    output DATA_O33;
    output DATA_O34;
    output DATA_O35;
    output DATA_O36;
    output DATA_O37;
    output DATA_O38;
    output DATA_O39;
    output DATA_O4;
    output DATA_O40;
    output DATA_O41;
    output DATA_O42;
    output DATA_O43;
    output DATA_O44;
    output DATA_O45;
    output DATA_O46;
    output DATA_O47;
    output DATA_O48;
    output DATA_O49;
    output DATA_O5;
    output DATA_O50;
    output DATA_O51;
    output DATA_O52;
    output DATA_O53;
    output DATA_O54;
    output DATA_O55;
    output DATA_O56;
    output DATA_O57;
    output DATA_O58;
    output DATA_O59;
    output DATA_O6;
    output DATA_O60;
    output DATA_O61;
    output DATA_O62;
    output DATA_O63;
    output DATA_O64;
    output DATA_O7;
    output DATA_O8;
    output DATA_O9;
    input DEC_E_I;
    input DSCR_E_I;
    output D_ERR_O1;
    output D_ERR_O2;
    output D_ERR_O3;
    output D_ERR_O4;
    output D_ERR_O5;
    output D_ERR_O6;
    output D_ERR_O7;
    output D_ERR_O8;
    inout [9:0] LINK;
    output LOCK_O;
    output LOS_O;
    output NIT_O1;
    output NIT_O2;
    output NIT_O3;
    output NIT_O4;
    output NIT_O5;
    output NIT_O6;
    output NIT_O7;
    output NIT_O8;
    input OVS_BS_I1;
    input OVS_BS_I2;
    input PLL_RN_I;
    input REP_E_I;
    input RST_N_I;
    input RX_I;
    input TST_I1;
    input TST_I2;
    input TST_I3;
    input TST_I4;
    output TST_O1;
    output TST_O2;
    output TST_O3;
    output TST_O4;
    output TST_O5;
    output TST_O6;
    output TST_O7;
    output TST_O8;
    parameter location = "";
    parameter pcs_8b_dscr_sel = 1'b0;
    parameter pcs_align_bypass = 1'b0;
    parameter pcs_buffers_bypass = 1'b0;
    parameter pcs_buffers_use_cdc = 1'b0;
    parameter pcs_bypass_pma_cdc = 1'b0;
    parameter pcs_bypass_usr_cdc = 1'b0;
    parameter pcs_comma_mask = 10'b0000000000;
    parameter pcs_debug_en = 1'b0;
    parameter pcs_dec_bypass = 1'b0;
    parameter pcs_dscr_bypass = 1'b0;
    parameter pcs_el_buff_diff_bef_comp = 3'b000;
    parameter pcs_el_buff_max_comp = 3'b000;
    parameter pcs_el_buff_only_one_skp = 1'b0;
    parameter pcs_el_buff_skp_char_0 = 9'b000000000;
    parameter pcs_el_buff_skp_char_1 = 9'b000000000;
    parameter pcs_el_buff_skp_char_2 = 9'b000000000;
    parameter pcs_el_buff_skp_char_3 = 9'b000000000;
    parameter pcs_el_buff_skp_header_0 = 9'b000000000;
    parameter pcs_el_buff_skp_header_1 = 9'b000000000;
    parameter pcs_el_buff_skp_header_2 = 9'b000000000;
    parameter pcs_el_buff_skp_header_3 = 9'b000000000;
    parameter pcs_el_buff_skp_header_size = 2'b00;
    parameter pcs_el_buff_skp_seq_size = 2'b00;
    parameter pcs_el_buff_underflow_handle = 1'b0;
    parameter pcs_fsm_sel = 2'b00;
    parameter pcs_fsm_watchdog_en = 1'b0;
    parameter pcs_loopback = 1'b0;
    parameter pcs_m_comma_en = 1'b0;
    parameter pcs_m_comma_val = 10'b0000000000;
    parameter pcs_nb_comma_bef_realign = 2'b00;
    parameter pcs_p_comma_en = 1'b0;
    parameter pcs_p_comma_val = 10'b0000000000;
    parameter pcs_polarity = 1'b0;
    parameter pcs_protocol_size = 1'b0;
    parameter pcs_replace_bypass = 1'b0;
    parameter pcs_sync_supported = 1'b0;
    parameter pma_cdr_cp = 4'b0000;
    parameter pma_clk_pos = 1'b0;
    parameter pma_ctrl_term = 6'b000000;
    parameter pma_loopback = 1'b0;
    parameter pma_pll_cpump_n = 3'b000;
    parameter pma_pll_divf = 2'b00;
    parameter pma_pll_divf_en_n = 1'b0;
    parameter pma_pll_divm = 2'b00;
    parameter pma_pll_divm_en_n = 1'b0;
    parameter pma_pll_divn = 1'b0;
    parameter pma_pll_divn_en_n = 1'b0;
    parameter test = 2'b00;
endmodule

(* blackbox *)
module NX_CRX_U(DSCR_E_I, DEC_E_I, ALIGN_E_I, ALIGN_S_I, REP_E_I, BUF_R_I, OVS_BS_I1, OVS_BS_I2, RST_N_I, PMA_RSTN_I, MEYE_RST_I, PWDN_N_I, DBG_S_I1, DBG_S_I2, DBG_S_I3, DATA_O1, DATA_O2, DATA_O3, DATA_O4, DATA_O5, DATA_O6
, DATA_O7, DATA_O8, DATA_O9, DATA_O10, DATA_O11, DATA_O12, DATA_O13, DATA_O14, DATA_O15, DATA_O16, DATA_O17, DATA_O18, DATA_O19, DATA_O20, DATA_O21, DATA_O22, DATA_O23, DATA_O24, DATA_O25, DATA_O26, DATA_O27
, DATA_O28, DATA_O29, DATA_O30, DATA_O31, DATA_O32, DATA_O33, DATA_O34, DATA_O35, DATA_O36, DATA_O37, DATA_O38, DATA_O39, DATA_O40, DATA_O41, DATA_O42, DATA_O43, DATA_O44, DATA_O45, DATA_O46, DATA_O47, DATA_O48
, DATA_O49, DATA_O50, DATA_O51, DATA_O52, DATA_O53, DATA_O54, DATA_O55, DATA_O56, DATA_O57, DATA_O58, DATA_O59, DATA_O60, DATA_O61, DATA_O62, DATA_O63, DATA_O64, CH_COM_O1, CH_COM_O2, CH_COM_O3, CH_COM_O4, CH_COM_O5
, CH_COM_O6, CH_COM_O7, CH_COM_O8, CH_K_O1, CH_K_O2, CH_K_O3, CH_K_O4, CH_K_O5, CH_K_O6, CH_K_O7, CH_K_O8, NIT_O1, NIT_O2, NIT_O3, NIT_O4, NIT_O5, NIT_O6, NIT_O7, NIT_O8, D_ERR_O1, D_ERR_O2
, D_ERR_O3, D_ERR_O4, D_ERR_O5, D_ERR_O6, D_ERR_O7, D_ERR_O8, CH_A_O1, CH_A_O2, CH_A_O3, CH_A_O4, CH_A_O5, CH_A_O6, CH_A_O7, CH_A_O8, CH_F_O1, CH_F_O2, CH_F_O3, CH_F_O4, CH_F_O5, CH_F_O6, CH_F_O7
, CH_F_O8, ALIGN_O, VREALIGN_O, BUSY_O, TST_O1, TST_O2, TST_O3, TST_O4, TST_O5, TST_O6, TST_O7, TST_O8, LOS_O, LL_FLOCK_O, LL_SLOCK_O, PLL_LOCK_O, PLL_LOCKT_O, LINK);
    input ALIGN_E_I;
    output ALIGN_O;
    input ALIGN_S_I;
    input BUF_R_I;
    output BUSY_O;
    output CH_A_O1;
    output CH_A_O2;
    output CH_A_O3;
    output CH_A_O4;
    output CH_A_O5;
    output CH_A_O6;
    output CH_A_O7;
    output CH_A_O8;
    output CH_COM_O1;
    output CH_COM_O2;
    output CH_COM_O3;
    output CH_COM_O4;
    output CH_COM_O5;
    output CH_COM_O6;
    output CH_COM_O7;
    output CH_COM_O8;
    output CH_F_O1;
    output CH_F_O2;
    output CH_F_O3;
    output CH_F_O4;
    output CH_F_O5;
    output CH_F_O6;
    output CH_F_O7;
    output CH_F_O8;
    output CH_K_O1;
    output CH_K_O2;
    output CH_K_O3;
    output CH_K_O4;
    output CH_K_O5;
    output CH_K_O6;
    output CH_K_O7;
    output CH_K_O8;
    output DATA_O1;
    output DATA_O10;
    output DATA_O11;
    output DATA_O12;
    output DATA_O13;
    output DATA_O14;
    output DATA_O15;
    output DATA_O16;
    output DATA_O17;
    output DATA_O18;
    output DATA_O19;
    output DATA_O2;
    output DATA_O20;
    output DATA_O21;
    output DATA_O22;
    output DATA_O23;
    output DATA_O24;
    output DATA_O25;
    output DATA_O26;
    output DATA_O27;
    output DATA_O28;
    output DATA_O29;
    output DATA_O3;
    output DATA_O30;
    output DATA_O31;
    output DATA_O32;
    output DATA_O33;
    output DATA_O34;
    output DATA_O35;
    output DATA_O36;
    output DATA_O37;
    output DATA_O38;
    output DATA_O39;
    output DATA_O4;
    output DATA_O40;
    output DATA_O41;
    output DATA_O42;
    output DATA_O43;
    output DATA_O44;
    output DATA_O45;
    output DATA_O46;
    output DATA_O47;
    output DATA_O48;
    output DATA_O49;
    output DATA_O5;
    output DATA_O50;
    output DATA_O51;
    output DATA_O52;
    output DATA_O53;
    output DATA_O54;
    output DATA_O55;
    output DATA_O56;
    output DATA_O57;
    output DATA_O58;
    output DATA_O59;
    output DATA_O6;
    output DATA_O60;
    output DATA_O61;
    output DATA_O62;
    output DATA_O63;
    output DATA_O64;
    output DATA_O7;
    output DATA_O8;
    output DATA_O9;
    input DBG_S_I1;
    input DBG_S_I2;
    input DBG_S_I3;
    input DEC_E_I;
    input DSCR_E_I;
    output D_ERR_O1;
    output D_ERR_O2;
    output D_ERR_O3;
    output D_ERR_O4;
    output D_ERR_O5;
    output D_ERR_O6;
    output D_ERR_O7;
    output D_ERR_O8;
    inout [9:0] LINK;
    output LL_FLOCK_O;
    output LL_SLOCK_O;
    output LOS_O;
    input MEYE_RST_I;
    output NIT_O1;
    output NIT_O2;
    output NIT_O3;
    output NIT_O4;
    output NIT_O5;
    output NIT_O6;
    output NIT_O7;
    output NIT_O8;
    input OVS_BS_I1;
    input OVS_BS_I2;
    output PLL_LOCKT_O;
    output PLL_LOCK_O;
    input PMA_RSTN_I;
    input PWDN_N_I;
    input REP_E_I;
    input RST_N_I;
    output TST_O1;
    output TST_O2;
    output TST_O3;
    output TST_O4;
    output TST_O5;
    output TST_O6;
    output TST_O7;
    output TST_O8;
    output VREALIGN_O;
    parameter gearbox_en = 1'b0;
    parameter gearbox_mode = 1'b0;
    parameter location = "";
    parameter pcs_8b_dscr_sel = 1'b0;
    parameter pcs_align_bypass = 1'b0;
    parameter pcs_buffers_bypass = 1'b0;
    parameter pcs_buffers_use_cdc = 1'b0;
    parameter pcs_bypass_pma_cdc = 1'b0;
    parameter pcs_bypass_usr_cdc = 1'b0;
    parameter pcs_comma_mask = 10'b0000000000;
    parameter pcs_debug_en = 1'b0;
    parameter pcs_dec_bypass = 1'b0;
    parameter pcs_dscr_bypass = 1'b0;
    parameter pcs_el_buff_diff_bef_comp = 4'b0000;
    parameter pcs_el_buff_max_comp = 4'b0000;
    parameter pcs_el_buff_only_one_skp = 1'b0;
    parameter pcs_el_buff_skp_char_0 = 9'b000000000;
    parameter pcs_el_buff_skp_char_1 = 9'b000000000;
    parameter pcs_el_buff_skp_char_2 = 9'b000000000;
    parameter pcs_el_buff_skp_char_3 = 9'b000000000;
    parameter pcs_el_buff_skp_header_0 = 9'b000000000;
    parameter pcs_el_buff_skp_header_1 = 9'b000000000;
    parameter pcs_el_buff_skp_header_2 = 9'b000000000;
    parameter pcs_el_buff_skp_header_3 = 9'b000000000;
    parameter pcs_el_buff_skp_header_size = 2'b00;
    parameter pcs_el_buff_skp_seq_size = 2'b00;
    parameter pcs_fsm_sel = 2'b00;
    parameter pcs_fsm_watchdog_en = 1'b0;
    parameter pcs_loopback = 1'b0;
    parameter pcs_m_comma_en = 1'b0;
    parameter pcs_m_comma_val = 10'b0000000000;
    parameter pcs_nb_comma_bef_realign = 2'b00;
    parameter pcs_p_comma_en = 1'b0;
    parameter pcs_p_comma_val = 10'b0000000000;
    parameter pcs_polarity = 1'b0;
    parameter pcs_protocol_size = 1'b0;
    parameter pcs_replace_bypass = 1'b0;
    parameter pcs_sync_supported = 1'b0;
    parameter pma_cdr_cp = 4'b0000;
    parameter pma_clk_pos = 1'b0;
    parameter pma_coarse_ppm = 3'b000;
    parameter pma_ctrl_term = 6'b000000;
    parameter pma_dco_divl = 2'b00;
    parameter pma_dco_divm = 1'b0;
    parameter pma_dco_divn = 2'b00;
    parameter pma_dco_reg_res = 2'b00;
    parameter pma_dco_vref_sel = 1'b0;
    parameter pma_fine_ppm = 3'b000;
    parameter pma_loopback = 1'b0;
    parameter pma_m_eye_ppm = 3'b000;
    parameter pma_peak_detect_cmd = 2'b00;
    parameter pma_peak_detect_on = 1'b0;
    parameter pma_pll_cpump_n = 3'b000;
    parameter pma_pll_divf = 2'b00;
    parameter pma_pll_divf_en_n = 1'b0;
    parameter pma_pll_divm = 2'b00;
    parameter pma_pll_divm_en_n = 1'b0;
    parameter pma_pll_divn = 1'b0;
    parameter pma_pll_divn_en_n = 1'b0;
endmodule

(* blackbox *)
module NX_CTX_L(ENC_E_I1, ENC_E_I2, ENC_E_I3, ENC_E_I4, ENC_E_I5, ENC_E_I6, ENC_E_I7, ENC_E_I8, CH_K_I1, CH_K_I2, CH_K_I3, CH_K_I4, CH_K_I5, CH_K_I6, CH_K_I7, CH_K_I8, SCR_E_I1, SCR_E_I2, SCR_E_I3, SCR_E_I4, SCR_E_I5
, SCR_E_I6, SCR_E_I7, SCR_E_I8, EOMF_I1, EOMF_I2, EOMF_I3, EOMF_I4, EOMF_I5, EOMF_I6, EOMF_I7, EOMF_I8, EOF_I1, EOF_I2, EOF_I3, EOF_I4, EOF_I5, EOF_I6, EOF_I7, EOF_I8, REP_E_I, RST_N_I
, TST_I1, TST_I2, TST_I3, TST_I4, DATA_I1, DATA_I2, DATA_I3, DATA_I4, DATA_I5, DATA_I6, DATA_I7, DATA_I8, DATA_I9, DATA_I10, DATA_I11, DATA_I12, DATA_I13, DATA_I14, DATA_I15, DATA_I16, DATA_I17
, DATA_I18, DATA_I19, DATA_I20, DATA_I21, DATA_I22, DATA_I23, DATA_I24, DATA_I25, DATA_I26, DATA_I27, DATA_I28, DATA_I29, DATA_I30, DATA_I31, DATA_I32, DATA_I33, DATA_I34, DATA_I35, DATA_I36, DATA_I37, DATA_I38
, DATA_I39, DATA_I40, DATA_I41, DATA_I42, DATA_I43, DATA_I44, DATA_I45, DATA_I46, DATA_I47, DATA_I48, DATA_I49, DATA_I50, DATA_I51, DATA_I52, DATA_I53, DATA_I54, DATA_I55, DATA_I56, DATA_I57, DATA_I58, DATA_I59
, DATA_I60, DATA_I61, DATA_I62, DATA_I63, DATA_I64, TST_O1, TST_O2, TST_O3, TST_O4, BUSY_O, CLK_E_I, TX_O, LINK);
    output BUSY_O;
    input CH_K_I1;
    input CH_K_I2;
    input CH_K_I3;
    input CH_K_I4;
    input CH_K_I5;
    input CH_K_I6;
    input CH_K_I7;
    input CH_K_I8;
    input CLK_E_I;
    input DATA_I1;
    input DATA_I10;
    input DATA_I11;
    input DATA_I12;
    input DATA_I13;
    input DATA_I14;
    input DATA_I15;
    input DATA_I16;
    input DATA_I17;
    input DATA_I18;
    input DATA_I19;
    input DATA_I2;
    input DATA_I20;
    input DATA_I21;
    input DATA_I22;
    input DATA_I23;
    input DATA_I24;
    input DATA_I25;
    input DATA_I26;
    input DATA_I27;
    input DATA_I28;
    input DATA_I29;
    input DATA_I3;
    input DATA_I30;
    input DATA_I31;
    input DATA_I32;
    input DATA_I33;
    input DATA_I34;
    input DATA_I35;
    input DATA_I36;
    input DATA_I37;
    input DATA_I38;
    input DATA_I39;
    input DATA_I4;
    input DATA_I40;
    input DATA_I41;
    input DATA_I42;
    input DATA_I43;
    input DATA_I44;
    input DATA_I45;
    input DATA_I46;
    input DATA_I47;
    input DATA_I48;
    input DATA_I49;
    input DATA_I5;
    input DATA_I50;
    input DATA_I51;
    input DATA_I52;
    input DATA_I53;
    input DATA_I54;
    input DATA_I55;
    input DATA_I56;
    input DATA_I57;
    input DATA_I58;
    input DATA_I59;
    input DATA_I6;
    input DATA_I60;
    input DATA_I61;
    input DATA_I62;
    input DATA_I63;
    input DATA_I64;
    input DATA_I7;
    input DATA_I8;
    input DATA_I9;
    input ENC_E_I1;
    input ENC_E_I2;
    input ENC_E_I3;
    input ENC_E_I4;
    input ENC_E_I5;
    input ENC_E_I6;
    input ENC_E_I7;
    input ENC_E_I8;
    input EOF_I1;
    input EOF_I2;
    input EOF_I3;
    input EOF_I4;
    input EOF_I5;
    input EOF_I6;
    input EOF_I7;
    input EOF_I8;
    input EOMF_I1;
    input EOMF_I2;
    input EOMF_I3;
    input EOMF_I4;
    input EOMF_I5;
    input EOMF_I6;
    input EOMF_I7;
    input EOMF_I8;
    inout [19:0] LINK;
    input REP_E_I;
    input RST_N_I;
    input SCR_E_I1;
    input SCR_E_I2;
    input SCR_E_I3;
    input SCR_E_I4;
    input SCR_E_I5;
    input SCR_E_I6;
    input SCR_E_I7;
    input SCR_E_I8;
    input TST_I1;
    input TST_I2;
    input TST_I3;
    input TST_I4;
    output TST_O1;
    output TST_O2;
    output TST_O3;
    output TST_O4;
    output TX_O;
    parameter location = "";
    parameter pcs_8b_scr_sel = 1'b0;
    parameter pcs_bypass_pma_cdc = 1'b0;
    parameter pcs_bypass_usr_cdc = 1'b0;
    parameter pcs_enc_bypass = 1'b0;
    parameter pcs_esistream_fsm_en = 1'b0;
    parameter pcs_loopback = 1'b0;
    parameter pcs_polarity = 1'b0;
    parameter pcs_protocol_size = 1'b0;
    parameter pcs_replace_bypass = 1'b0;
    parameter pcs_scr_bypass = 1'b0;
    parameter pcs_scr_init = 17'b00000000000000000;
    parameter pcs_sync_supported = 1'b0;
    parameter pma_clk_pos = 1'b0;
    parameter pma_loopback = 1'b0;
    parameter test = 2'b00;
endmodule

(* blackbox *)
module NX_CTX_U(ENC_E_I1, ENC_E_I2, ENC_E_I3, ENC_E_I4, ENC_E_I5, ENC_E_I6, ENC_E_I7, ENC_E_I8, CH_K_I1, CH_K_I2, CH_K_I3, CH_K_I4, CH_K_I5, CH_K_I6, CH_K_I7, CH_K_I8, SCR_E_I1, SCR_E_I2, SCR_E_I3, SCR_E_I4, SCR_E_I5
, SCR_E_I6, SCR_E_I7, SCR_E_I8, EOMF_I1, EOMF_I2, EOMF_I3, EOMF_I4, EOMF_I5, EOMF_I6, EOMF_I7, EOMF_I8, EOF_I1, EOF_I2, EOF_I3, EOF_I4, EOF_I5, EOF_I6, EOF_I7, EOF_I8, REP_E_I, RST_N_I
, DATA_I1, DATA_I2, DATA_I3, DATA_I4, DATA_I5, DATA_I6, DATA_I7, DATA_I8, DATA_I9, DATA_I10, DATA_I11, DATA_I12, DATA_I13, DATA_I14, DATA_I15, DATA_I16, DATA_I17, DATA_I18, DATA_I19, DATA_I20, DATA_I21
, DATA_I22, DATA_I23, DATA_I24, DATA_I25, DATA_I26, DATA_I27, DATA_I28, DATA_I29, DATA_I30, DATA_I31, DATA_I32, DATA_I33, DATA_I34, DATA_I35, DATA_I36, DATA_I37, DATA_I38, DATA_I39, DATA_I40, DATA_I41, DATA_I42
, DATA_I43, DATA_I44, DATA_I45, DATA_I46, DATA_I47, DATA_I48, DATA_I49, DATA_I50, DATA_I51, DATA_I52, DATA_I53, DATA_I54, DATA_I55, DATA_I56, DATA_I57, DATA_I58, DATA_I59, DATA_I60, DATA_I61, DATA_I62, DATA_I63
, DATA_I64, BUSY_O, INV_K_O, PWDN_N_I, CLK_E_I, CLK_O, LINK);
    output BUSY_O;
    input CH_K_I1;
    input CH_K_I2;
    input CH_K_I3;
    input CH_K_I4;
    input CH_K_I5;
    input CH_K_I6;
    input CH_K_I7;
    input CH_K_I8;
    input CLK_E_I;
    output CLK_O;
    input DATA_I1;
    input DATA_I10;
    input DATA_I11;
    input DATA_I12;
    input DATA_I13;
    input DATA_I14;
    input DATA_I15;
    input DATA_I16;
    input DATA_I17;
    input DATA_I18;
    input DATA_I19;
    input DATA_I2;
    input DATA_I20;
    input DATA_I21;
    input DATA_I22;
    input DATA_I23;
    input DATA_I24;
    input DATA_I25;
    input DATA_I26;
    input DATA_I27;
    input DATA_I28;
    input DATA_I29;
    input DATA_I3;
    input DATA_I30;
    input DATA_I31;
    input DATA_I32;
    input DATA_I33;
    input DATA_I34;
    input DATA_I35;
    input DATA_I36;
    input DATA_I37;
    input DATA_I38;
    input DATA_I39;
    input DATA_I4;
    input DATA_I40;
    input DATA_I41;
    input DATA_I42;
    input DATA_I43;
    input DATA_I44;
    input DATA_I45;
    input DATA_I46;
    input DATA_I47;
    input DATA_I48;
    input DATA_I49;
    input DATA_I5;
    input DATA_I50;
    input DATA_I51;
    input DATA_I52;
    input DATA_I53;
    input DATA_I54;
    input DATA_I55;
    input DATA_I56;
    input DATA_I57;
    input DATA_I58;
    input DATA_I59;
    input DATA_I6;
    input DATA_I60;
    input DATA_I61;
    input DATA_I62;
    input DATA_I63;
    input DATA_I64;
    input DATA_I7;
    input DATA_I8;
    input DATA_I9;
    input ENC_E_I1;
    input ENC_E_I2;
    input ENC_E_I3;
    input ENC_E_I4;
    input ENC_E_I5;
    input ENC_E_I6;
    input ENC_E_I7;
    input ENC_E_I8;
    input EOF_I1;
    input EOF_I2;
    input EOF_I3;
    input EOF_I4;
    input EOF_I5;
    input EOF_I6;
    input EOF_I7;
    input EOF_I8;
    input EOMF_I1;
    input EOMF_I2;
    input EOMF_I3;
    input EOMF_I4;
    input EOMF_I5;
    input EOMF_I6;
    input EOMF_I7;
    input EOMF_I8;
    output INV_K_O;
    inout [19:0] LINK;
    input PWDN_N_I;
    input REP_E_I;
    input RST_N_I;
    input SCR_E_I1;
    input SCR_E_I2;
    input SCR_E_I3;
    input SCR_E_I4;
    input SCR_E_I5;
    input SCR_E_I6;
    input SCR_E_I7;
    input SCR_E_I8;
    parameter gearbox_en = 1'b0;
    parameter gearbox_mode = 1'b0;
    parameter location = "";
    parameter pcs_8b_scr_sel = 1'b0;
    parameter pcs_bypass_pma_cdc = 1'b0;
    parameter pcs_bypass_usr_cdc = 1'b0;
    parameter pcs_enc_bypass = 1'b0;
    parameter pcs_esistream_fsm_en = 1'b0;
    parameter pcs_loopback = 1'b0;
    parameter pcs_polarity = 1'b0;
    parameter pcs_protocol_size = 1'b0;
    parameter pcs_replace_bypass = 1'b0;
    parameter pcs_scr_bypass = 1'b0;
    parameter pcs_scr_init = 17'b00000000000000000;
    parameter pcs_sync_supported = 1'b0;
    parameter pma_clk_pos = 1'b0;
    parameter pma_loopback = 1'b0;
endmodule

//(* blackbox *)
//module NX_CY(A1, A2, A3, A4, B1, B2, B3, B4, CI, CO, S1, S2, S3, S4);
//    input A1;
//    input A2;
//    input A3;
//    input A4;
//    input B1;
//    input B2;
//    input B3;
//    input B4;
//    input CI;
//    output CO;
//    output S1;
//    output S2;
//    output S3;
//    output S4;
//    parameter add_carry = 0;
//endmodule

(* blackbox *)
module NX_DES(FCK, SCK, R, IO, DCK, DRL, DIG, FZ, FLD, FLG, O, DS, DRA, DRI, DRO, DID);
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    input FCK;
    output FLD;
    output FLG;
    input FZ;
    input IO;
    output [4:0] O;
    input R;
    input SCK;
    parameter data_size = 5;
    parameter differential = "";
    parameter dpath_dynamic = 1'b0;
    parameter drive = "";
    parameter inputDelayLine = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

//(* blackbox *)
//module NX_DFF(I, CK, L, R, O);
//    input CK;
//    input I;
//    input L;
//    output O;
//    input R;
//    parameter dff_ctxt = 1'b0;
//    parameter dff_edge = 1'b0;
//    parameter dff_init = 1'b0;
//    parameter dff_load = 1'b0;
//    parameter dff_sync = 1'b0;
//    parameter dff_type = 1'b0;
//endmodule

(* blackbox *)
module NX_DFR(I, CK, L, R, O);
    input CK;
    input I;
    input L;
    output O;
    input R;
    parameter data_inv = 1'b0;
    parameter dff_edge = 1'b0;
    parameter dff_init = 1'b0;
    parameter dff_load = 1'b0;
    parameter dff_sync = 1'b0;
    parameter dff_type = 1'b0;
    parameter iobname = "";
    parameter location = "";
    parameter mode = 0;
    parameter path = 0;
    parameter ring = 0;
endmodule

(* blackbox *)
module NX_DSP(A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17, A18, A19, A20, A21
, A22, A23, A24, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15, B16, B17, B18
, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16, C17, C18, C19, C20, C21
, C22, C23, C24, C25, C26, C27, C28, C29, C30, C31, C32, C33, C34, C35, C36, CAI1, CAI2, CAI3, CAI4, CAI5, CAI6
, CAI7, CAI8, CAI9, CAI10, CAI11, CAI12, CAI13, CAI14, CAI15, CAI16, CAI17, CAI18, CAO1, CAO2, CAO3, CAO4, CAO5, CAO6, CAO7, CAO8, CAO9
, CAO10, CAO11, CAO12, CAO13, CAO14, CAO15, CAO16, CAO17, CAO18, CBI1, CBI2, CBI3, CBI4, CBI5, CBI6, CBI7, CBI8, CBI9, CBI10, CBI11, CBI12
, CBI13, CBI14, CBI15, CBI16, CBI17, CBI18, CBO1, CBO2, CBO3, CBO4, CBO5, CBO6, CBO7, CBO8, CBO9, CBO10, CBO11, CBO12, CBO13, CBO14, CBO15
, CBO16, CBO17, CBO18, CCI, CCO, CI, CK, CO, CO37, CO49, CZI1, CZI2, CZI3, CZI4, CZI5, CZI6, CZI7, CZI8, CZI9, CZI10, CZI11
, CZI12, CZI13, CZI14, CZI15, CZI16, CZI17, CZI18, CZI19, CZI20, CZI21, CZI22, CZI23, CZI24, CZI25, CZI26, CZI27, CZI28, CZI29, CZI30, CZI31, CZI32
, CZI33, CZI34, CZI35, CZI36, CZI37, CZI38, CZI39, CZI40, CZI41, CZI42, CZI43, CZI44, CZI45, CZI46, CZI47, CZI48, CZI49, CZI50, CZI51, CZI52, CZI53
, CZI54, CZI55, CZI56, CZO1, CZO2, CZO3, CZO4, CZO5, CZO6, CZO7, CZO8, CZO9, CZO10, CZO11, CZO12, CZO13, CZO14, CZO15, CZO16, CZO17, CZO18
, CZO19, CZO20, CZO21, CZO22, CZO23, CZO24, CZO25, CZO26, CZO27, CZO28, CZO29, CZO30, CZO31, CZO32, CZO33, CZO34, CZO35, CZO36, CZO37, CZO38, CZO39
, CZO40, CZO41, CZO42, CZO43, CZO44, CZO45, CZO46, CZO47, CZO48, CZO49, CZO50, CZO51, CZO52, CZO53, CZO54, CZO55, CZO56, D1, D2, D3, D4
, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, D16, D17, D18, OVF, R, RZ, WE, Z1, Z2, Z3
, Z4, Z5, Z6, Z7, Z8, Z9, Z10, Z11, Z12, Z13, Z14, Z15, Z16, Z17, Z18, Z19, Z20, Z21, Z22, Z23, Z24
, Z25, Z26, Z27, Z28, Z29, Z30, Z31, Z32, Z33, Z34, Z35, Z36, Z37, Z38, Z39, Z40, Z41, Z42, Z43, Z44, Z45
, Z46, Z47, Z48, Z49, Z50, Z51, Z52, Z53, Z54, Z55, Z56);
    input A1;
    input A10;
    input A11;
    input A12;
    input A13;
    input A14;
    input A15;
    input A16;
    input A17;
    input A18;
    input A19;
    input A2;
    input A20;
    input A21;
    input A22;
    input A23;
    input A24;
    input A3;
    input A4;
    input A5;
    input A6;
    input A7;
    input A8;
    input A9;
    input B1;
    input B10;
    input B11;
    input B12;
    input B13;
    input B14;
    input B15;
    input B16;
    input B17;
    input B18;
    input B2;
    input B3;
    input B4;
    input B5;
    input B6;
    input B7;
    input B8;
    input B9;
    input C1;
    input C10;
    input C11;
    input C12;
    input C13;
    input C14;
    input C15;
    input C16;
    input C17;
    input C18;
    input C19;
    input C2;
    input C20;
    input C21;
    input C22;
    input C23;
    input C24;
    input C25;
    input C26;
    input C27;
    input C28;
    input C29;
    input C3;
    input C30;
    input C31;
    input C32;
    input C33;
    input C34;
    input C35;
    input C36;
    input C4;
    input C5;
    input C6;
    input C7;
    input C8;
    input C9;
    input CAI1;
    input CAI10;
    input CAI11;
    input CAI12;
    input CAI13;
    input CAI14;
    input CAI15;
    input CAI16;
    input CAI17;
    input CAI18;
    input CAI2;
    input CAI3;
    input CAI4;
    input CAI5;
    input CAI6;
    input CAI7;
    input CAI8;
    input CAI9;
    output CAO1;
    output CAO10;
    output CAO11;
    output CAO12;
    output CAO13;
    output CAO14;
    output CAO15;
    output CAO16;
    output CAO17;
    output CAO18;
    output CAO2;
    output CAO3;
    output CAO4;
    output CAO5;
    output CAO6;
    output CAO7;
    output CAO8;
    output CAO9;
    input CBI1;
    input CBI10;
    input CBI11;
    input CBI12;
    input CBI13;
    input CBI14;
    input CBI15;
    input CBI16;
    input CBI17;
    input CBI18;
    input CBI2;
    input CBI3;
    input CBI4;
    input CBI5;
    input CBI6;
    input CBI7;
    input CBI8;
    input CBI9;
    output CBO1;
    output CBO10;
    output CBO11;
    output CBO12;
    output CBO13;
    output CBO14;
    output CBO15;
    output CBO16;
    output CBO17;
    output CBO18;
    output CBO2;
    output CBO3;
    output CBO4;
    output CBO5;
    output CBO6;
    output CBO7;
    output CBO8;
    output CBO9;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO;
    output CO37;
    output CO49;
    input CZI1;
    input CZI10;
    input CZI11;
    input CZI12;
    input CZI13;
    input CZI14;
    input CZI15;
    input CZI16;
    input CZI17;
    input CZI18;
    input CZI19;
    input CZI2;
    input CZI20;
    input CZI21;
    input CZI22;
    input CZI23;
    input CZI24;
    input CZI25;
    input CZI26;
    input CZI27;
    input CZI28;
    input CZI29;
    input CZI3;
    input CZI30;
    input CZI31;
    input CZI32;
    input CZI33;
    input CZI34;
    input CZI35;
    input CZI36;
    input CZI37;
    input CZI38;
    input CZI39;
    input CZI4;
    input CZI40;
    input CZI41;
    input CZI42;
    input CZI43;
    input CZI44;
    input CZI45;
    input CZI46;
    input CZI47;
    input CZI48;
    input CZI49;
    input CZI5;
    input CZI50;
    input CZI51;
    input CZI52;
    input CZI53;
    input CZI54;
    input CZI55;
    input CZI56;
    input CZI6;
    input CZI7;
    input CZI8;
    input CZI9;
    output CZO1;
    output CZO10;
    output CZO11;
    output CZO12;
    output CZO13;
    output CZO14;
    output CZO15;
    output CZO16;
    output CZO17;
    output CZO18;
    output CZO19;
    output CZO2;
    output CZO20;
    output CZO21;
    output CZO22;
    output CZO23;
    output CZO24;
    output CZO25;
    output CZO26;
    output CZO27;
    output CZO28;
    output CZO29;
    output CZO3;
    output CZO30;
    output CZO31;
    output CZO32;
    output CZO33;
    output CZO34;
    output CZO35;
    output CZO36;
    output CZO37;
    output CZO38;
    output CZO39;
    output CZO4;
    output CZO40;
    output CZO41;
    output CZO42;
    output CZO43;
    output CZO44;
    output CZO45;
    output CZO46;
    output CZO47;
    output CZO48;
    output CZO49;
    output CZO5;
    output CZO50;
    output CZO51;
    output CZO52;
    output CZO53;
    output CZO54;
    output CZO55;
    output CZO56;
    output CZO6;
    output CZO7;
    output CZO8;
    output CZO9;
    input D1;
    input D10;
    input D11;
    input D12;
    input D13;
    input D14;
    input D15;
    input D16;
    input D17;
    input D18;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input D8;
    input D9;
    output OVF;
    input R;
    input RZ;
    input WE;
    output Z1;
    output Z10;
    output Z11;
    output Z12;
    output Z13;
    output Z14;
    output Z15;
    output Z16;
    output Z17;
    output Z18;
    output Z19;
    output Z2;
    output Z20;
    output Z21;
    output Z22;
    output Z23;
    output Z24;
    output Z25;
    output Z26;
    output Z27;
    output Z28;
    output Z29;
    output Z3;
    output Z30;
    output Z31;
    output Z32;
    output Z33;
    output Z34;
    output Z35;
    output Z36;
    output Z37;
    output Z38;
    output Z39;
    output Z4;
    output Z40;
    output Z41;
    output Z42;
    output Z43;
    output Z44;
    output Z45;
    output Z46;
    output Z47;
    output Z48;
    output Z49;
    output Z5;
    output Z50;
    output Z51;
    output Z52;
    output Z53;
    output Z54;
    output Z55;
    output Z56;
    output Z6;
    output Z7;
    output Z8;
    output Z9;
    parameter raw_config0 = 20'b00000000000000000000;
    parameter raw_config1 = 19'b0000000000000000000;
    parameter raw_config2 = 13'b0000000000000;
    parameter raw_config3 = 7'b0000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_DSP_L(A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17, A18, A19, A20, A21
, A22, A23, A24, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15, B16, B17, B18
, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16, C17, C18, C19, C20, C21
, C22, C23, C24, C25, C26, C27, C28, C29, C30, C31, C32, C33, C34, C35, C36, CAI1, CAI2, CAI3, CAI4, CAI5, CAI6
, CAI7, CAI8, CAI9, CAI10, CAI11, CAI12, CAI13, CAI14, CAI15, CAI16, CAI17, CAI18, CAI19, CAI20, CAI21, CAI22, CAI23, CAI24, CAO1, CAO2, CAO3
, CAO4, CAO5, CAO6, CAO7, CAO8, CAO9, CAO10, CAO11, CAO12, CAO13, CAO14, CAO15, CAO16, CAO17, CAO18, CAO19, CAO20, CAO21, CAO22, CAO23, CAO24
, CBI1, CBI2, CBI3, CBI4, CBI5, CBI6, CBI7, CBI8, CBI9, CBI10, CBI11, CBI12, CBI13, CBI14, CBI15, CBI16, CBI17, CBI18, CBO1, CBO2, CBO3
, CBO4, CBO5, CBO6, CBO7, CBO8, CBO9, CBO10, CBO11, CBO12, CBO13, CBO14, CBO15, CBO16, CBO17, CBO18, CCI, CCO, CI, CK, CO, CO37
, CO57, CZI1, CZI2, CZI3, CZI4, CZI5, CZI6, CZI7, CZI8, CZI9, CZI10, CZI11, CZI12, CZI13, CZI14, CZI15, CZI16, CZI17, CZI18, CZI19, CZI20
, CZI21, CZI22, CZI23, CZI24, CZI25, CZI26, CZI27, CZI28, CZI29, CZI30, CZI31, CZI32, CZI33, CZI34, CZI35, CZI36, CZI37, CZI38, CZI39, CZI40, CZI41
, CZI42, CZI43, CZI44, CZI45, CZI46, CZI47, CZI48, CZI49, CZI50, CZI51, CZI52, CZI53, CZI54, CZI55, CZI56, CZO1, CZO2, CZO3, CZO4, CZO5, CZO6
, CZO7, CZO8, CZO9, CZO10, CZO11, CZO12, CZO13, CZO14, CZO15, CZO16, CZO17, CZO18, CZO19, CZO20, CZO21, CZO22, CZO23, CZO24, CZO25, CZO26, CZO27
, CZO28, CZO29, CZO30, CZO31, CZO32, CZO33, CZO34, CZO35, CZO36, CZO37, CZO38, CZO39, CZO40, CZO41, CZO42, CZO43, CZO44, CZO45, CZO46, CZO47, CZO48
, CZO49, CZO50, CZO51, CZO52, CZO53, CZO54, CZO55, CZO56, D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13
, D14, D15, D16, D17, D18, OVF, R, RZ, WE, Z1, Z2, Z3, Z4, Z5, Z6, Z7, Z8, Z9, Z10, Z11, Z12
, Z13, Z14, Z15, Z16, Z17, Z18, Z19, Z20, Z21, Z22, Z23, Z24, Z25, Z26, Z27, Z28, Z29, Z30, Z31, Z32, Z33
, Z34, Z35, Z36, Z37, Z38, Z39, Z40, Z41, Z42, Z43, Z44, Z45, Z46, Z47, Z48, Z49, Z50, Z51, Z52, Z53, Z54
, Z55, Z56);
    input A1;
    input A10;
    input A11;
    input A12;
    input A13;
    input A14;
    input A15;
    input A16;
    input A17;
    input A18;
    input A19;
    input A2;
    input A20;
    input A21;
    input A22;
    input A23;
    input A24;
    input A3;
    input A4;
    input A5;
    input A6;
    input A7;
    input A8;
    input A9;
    input B1;
    input B10;
    input B11;
    input B12;
    input B13;
    input B14;
    input B15;
    input B16;
    input B17;
    input B18;
    input B2;
    input B3;
    input B4;
    input B5;
    input B6;
    input B7;
    input B8;
    input B9;
    input C1;
    input C10;
    input C11;
    input C12;
    input C13;
    input C14;
    input C15;
    input C16;
    input C17;
    input C18;
    input C19;
    input C2;
    input C20;
    input C21;
    input C22;
    input C23;
    input C24;
    input C25;
    input C26;
    input C27;
    input C28;
    input C29;
    input C3;
    input C30;
    input C31;
    input C32;
    input C33;
    input C34;
    input C35;
    input C36;
    input C4;
    input C5;
    input C6;
    input C7;
    input C8;
    input C9;
    input CAI1;
    input CAI10;
    input CAI11;
    input CAI12;
    input CAI13;
    input CAI14;
    input CAI15;
    input CAI16;
    input CAI17;
    input CAI18;
    input CAI19;
    input CAI2;
    input CAI20;
    input CAI21;
    input CAI22;
    input CAI23;
    input CAI24;
    input CAI3;
    input CAI4;
    input CAI5;
    input CAI6;
    input CAI7;
    input CAI8;
    input CAI9;
    output CAO1;
    output CAO10;
    output CAO11;
    output CAO12;
    output CAO13;
    output CAO14;
    output CAO15;
    output CAO16;
    output CAO17;
    output CAO18;
    output CAO19;
    output CAO2;
    output CAO20;
    output CAO21;
    output CAO22;
    output CAO23;
    output CAO24;
    output CAO3;
    output CAO4;
    output CAO5;
    output CAO6;
    output CAO7;
    output CAO8;
    output CAO9;
    input CBI1;
    input CBI10;
    input CBI11;
    input CBI12;
    input CBI13;
    input CBI14;
    input CBI15;
    input CBI16;
    input CBI17;
    input CBI18;
    input CBI2;
    input CBI3;
    input CBI4;
    input CBI5;
    input CBI6;
    input CBI7;
    input CBI8;
    input CBI9;
    output CBO1;
    output CBO10;
    output CBO11;
    output CBO12;
    output CBO13;
    output CBO14;
    output CBO15;
    output CBO16;
    output CBO17;
    output CBO18;
    output CBO2;
    output CBO3;
    output CBO4;
    output CBO5;
    output CBO6;
    output CBO7;
    output CBO8;
    output CBO9;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO;
    output CO37;
    output CO57;
    input CZI1;
    input CZI10;
    input CZI11;
    input CZI12;
    input CZI13;
    input CZI14;
    input CZI15;
    input CZI16;
    input CZI17;
    input CZI18;
    input CZI19;
    input CZI2;
    input CZI20;
    input CZI21;
    input CZI22;
    input CZI23;
    input CZI24;
    input CZI25;
    input CZI26;
    input CZI27;
    input CZI28;
    input CZI29;
    input CZI3;
    input CZI30;
    input CZI31;
    input CZI32;
    input CZI33;
    input CZI34;
    input CZI35;
    input CZI36;
    input CZI37;
    input CZI38;
    input CZI39;
    input CZI4;
    input CZI40;
    input CZI41;
    input CZI42;
    input CZI43;
    input CZI44;
    input CZI45;
    input CZI46;
    input CZI47;
    input CZI48;
    input CZI49;
    input CZI5;
    input CZI50;
    input CZI51;
    input CZI52;
    input CZI53;
    input CZI54;
    input CZI55;
    input CZI56;
    input CZI6;
    input CZI7;
    input CZI8;
    input CZI9;
    output CZO1;
    output CZO10;
    output CZO11;
    output CZO12;
    output CZO13;
    output CZO14;
    output CZO15;
    output CZO16;
    output CZO17;
    output CZO18;
    output CZO19;
    output CZO2;
    output CZO20;
    output CZO21;
    output CZO22;
    output CZO23;
    output CZO24;
    output CZO25;
    output CZO26;
    output CZO27;
    output CZO28;
    output CZO29;
    output CZO3;
    output CZO30;
    output CZO31;
    output CZO32;
    output CZO33;
    output CZO34;
    output CZO35;
    output CZO36;
    output CZO37;
    output CZO38;
    output CZO39;
    output CZO4;
    output CZO40;
    output CZO41;
    output CZO42;
    output CZO43;
    output CZO44;
    output CZO45;
    output CZO46;
    output CZO47;
    output CZO48;
    output CZO49;
    output CZO5;
    output CZO50;
    output CZO51;
    output CZO52;
    output CZO53;
    output CZO54;
    output CZO55;
    output CZO56;
    output CZO6;
    output CZO7;
    output CZO8;
    output CZO9;
    input D1;
    input D10;
    input D11;
    input D12;
    input D13;
    input D14;
    input D15;
    input D16;
    input D17;
    input D18;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input D8;
    input D9;
    output OVF;
    input R;
    input RZ;
    input WE;
    output Z1;
    output Z10;
    output Z11;
    output Z12;
    output Z13;
    output Z14;
    output Z15;
    output Z16;
    output Z17;
    output Z18;
    output Z19;
    output Z2;
    output Z20;
    output Z21;
    output Z22;
    output Z23;
    output Z24;
    output Z25;
    output Z26;
    output Z27;
    output Z28;
    output Z29;
    output Z3;
    output Z30;
    output Z31;
    output Z32;
    output Z33;
    output Z34;
    output Z35;
    output Z36;
    output Z37;
    output Z38;
    output Z39;
    output Z4;
    output Z40;
    output Z41;
    output Z42;
    output Z43;
    output Z44;
    output Z45;
    output Z46;
    output Z47;
    output Z48;
    output Z49;
    output Z5;
    output Z50;
    output Z51;
    output Z52;
    output Z53;
    output Z54;
    output Z55;
    output Z56;
    output Z6;
    output Z7;
    output Z8;
    output Z9;
    parameter raw_config0 = 20'b00000000000000000000;
    parameter raw_config1 = 19'b0000000000000000000;
    parameter raw_config2 = 13'b0000000000000;
    parameter raw_config3 = 7'b0000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_DSP_L_SPLIT(CK, R, RZ, WE, CI, CCI, CO, CO36, CO56, OVF, CCO, A, B, C, D, Z, CAI, CBI, CZI, CAO, CBO
, CZO);
    input [23:0] A;
    input [17:0] B;
    input [35:0] C;
    input [23:0] CAI;
    output [23:0] CAO;
    input [17:0] CBI;
    output [17:0] CBO;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO;
    output CO36;
    output CO56;
    input [55:0] CZI;
    output [55:0] CZO;
    input [17:0] D;
    output OVF;
    input R;
    input RZ;
    input WE;
    output [55:0] Z;
    parameter ALU_DYNAMIC_OP = 1'b0;
    parameter ALU_MUX = 1'b0;
    parameter ALU_OP = 6'b000000;
    parameter CO_SEL = 1'b0;
    parameter ENABLE_PR_ALU_RST = 1'b0;
    parameter ENABLE_PR_A_RST = 1'b0;
    parameter ENABLE_PR_B_RST = 1'b0;
    parameter ENABLE_PR_CI_RST = 1'b0;
    parameter ENABLE_PR_CO_RST = 1'b0;
    parameter ENABLE_PR_C_RST = 1'b0;
    parameter ENABLE_PR_D_RST = 1'b0;
    parameter ENABLE_PR_MULT_RST = 1'b0;
    parameter ENABLE_PR_OV_RST = 1'b0;
    parameter ENABLE_PR_P_RST = 1'b0;
    parameter ENABLE_PR_X_RST = 1'b0;
    parameter ENABLE_PR_Y_RST = 1'b0;
    parameter ENABLE_PR_Z_RST = 1'b0;
    parameter ENABLE_SATURATION = 1'b0;
    parameter MUX_A = 1'b0;
    parameter MUX_B = 1'b0;
    parameter MUX_CI = 1'b0;
    parameter MUX_P = 1'b0;
    parameter MUX_X = 2'b00;
    parameter MUX_Y = 1'b0;
    parameter MUX_Z = 1'b0;
    parameter PRE_ADDER_OP = 1'b0;
    parameter PR_ALU_MUX = 1'b0;
    parameter PR_A_CASCADE_MUX = 2'b00;
    parameter PR_A_MUX = 2'b00;
    parameter PR_B_CASCADE_MUX = 2'b00;
    parameter PR_B_MUX = 2'b00;
    parameter PR_CI_MUX = 1'b0;
    parameter PR_CO_MUX = 1'b0;
    parameter PR_C_MUX = 1'b0;
    parameter PR_D_MUX = 1'b0;
    parameter PR_MULT_MUX = 1'b0;
    parameter PR_OV_MUX = 1'b0;
    parameter PR_P_MUX = 1'b0;
    parameter PR_X_MUX = 1'b0;
    parameter PR_Y_MUX = 1'b0;
    parameter PR_Z_MUX = 1'b0;
    parameter SATURATION_RANK = 6'b000000;
    parameter SIGNED_MODE = 1'b0;
    parameter Z_FEEDBACK_SHL12 = 1'b0;
endmodule

(* blackbox *)
module NX_DSP_L_WRAP(CCI, CCO, CI, CK, CO, CO37, CO57, OVF, R, RZ, WE, A, B, C, D, Z, CAI, CBI, CZI, CAO, CBO
, CZO);
    input [23:0] A;
    input [17:0] B;
    input [35:0] C;
    input [23:0] CAI;
    output [23:0] CAO;
    input [17:0] CBI;
    output [17:0] CBO;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO;
    output CO37;
    output CO57;
    input [55:0] CZI;
    output [55:0] CZO;
    input [17:0] D;
    output OVF;
    input R;
    input RZ;
    input WE;
    output [55:0] Z;
    parameter raw_config0 = 20'b00000000000000000000;
    parameter raw_config1 = 19'b0000000000000000000;
    parameter raw_config2 = 13'b0000000000000;
    parameter raw_config3 = 7'b0000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_DSP_SPLIT(CK, R, RZ, WE, CI, CCI, CO, CO36, CO48, OVF, CCO, A, B, C, D, Z, CAI, CBI, CZI, CAO, CBO
, CZO);
    input [23:0] A;
    input [17:0] B;
    input [35:0] C;
    input [17:0] CAI;
    output [17:0] CAO;
    input [17:0] CBI;
    output [17:0] CBO;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO;
    output CO36;
    output CO48;
    input [55:0] CZI;
    output [55:0] CZO;
    input [17:0] D;
    output OVF;
    input R;
    input RZ;
    input WE;
    output [55:0] Z;
    parameter ALU_DYNAMIC_OP = 1'b0;
    parameter ALU_MUX = 1'b0;
    parameter ALU_OP = 6'b000000;
    parameter CO_SEL = 1'b0;
    parameter ENABLE_PR_ALU_RST = 1'b0;
    parameter ENABLE_PR_A_RST = 1'b0;
    parameter ENABLE_PR_B_RST = 1'b0;
    parameter ENABLE_PR_CI_RST = 1'b0;
    parameter ENABLE_PR_CO_RST = 1'b0;
    parameter ENABLE_PR_C_RST = 1'b0;
    parameter ENABLE_PR_D_RST = 1'b0;
    parameter ENABLE_PR_MULT_RST = 1'b0;
    parameter ENABLE_PR_OV_RST = 1'b0;
    parameter ENABLE_PR_P_RST = 1'b0;
    parameter ENABLE_PR_X_RST = 1'b0;
    parameter ENABLE_PR_Y_RST = 1'b0;
    parameter ENABLE_PR_Z_RST = 1'b0;
    parameter ENABLE_SATURATION = 1'b0;
    parameter MUX_A = 1'b0;
    parameter MUX_B = 1'b0;
    parameter MUX_CI = 1'b0;
    parameter MUX_P = 1'b0;
    parameter MUX_X = 2'b00;
    parameter MUX_Y = 1'b0;
    parameter MUX_Z = 1'b0;
    parameter PRE_ADDER_OP = 1'b0;
    parameter PR_ALU_MUX = 1'b0;
    parameter PR_A_CASCADE_MUX = 2'b00;
    parameter PR_A_MUX = 2'b00;
    parameter PR_B_CASCADE_MUX = 2'b00;
    parameter PR_B_MUX = 2'b00;
    parameter PR_CI_MUX = 1'b0;
    parameter PR_CO_MUX = 1'b0;
    parameter PR_C_MUX = 1'b0;
    parameter PR_D_MUX = 1'b0;
    parameter PR_MULT_MUX = 1'b0;
    parameter PR_OV_MUX = 1'b0;
    parameter PR_P_MUX = 1'b0;
    parameter PR_X_MUX = 1'b0;
    parameter PR_Y_MUX = 1'b0;
    parameter PR_Z_MUX = 1'b0;
    parameter SATURATION_RANK = 6'b000000;
    parameter SIGNED_MODE = 1'b0;
    parameter Z_FEEDBACK_SHL12 = 1'b0;
endmodule

(* blackbox *)
module NX_DSP_U(A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17, A18, A19, A20, A21
, A22, A23, A24, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15, B16, B17, B18
, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16, C17, C18, C19, C20, C21
, C22, C23, C24, C25, C26, C27, C28, C29, C30, C31, C32, C33, C34, C35, C36, CAI1, CAI2, CAI3, CAI4, CAI5, CAI6
, CAI7, CAI8, CAI9, CAI10, CAI11, CAI12, CAI13, CAI14, CAI15, CAI16, CAI17, CAI18, CAI19, CAI20, CAI21, CAI22, CAI23, CAI24, CAO1, CAO2, CAO3
, CAO4, CAO5, CAO6, CAO7, CAO8, CAO9, CAO10, CAO11, CAO12, CAO13, CAO14, CAO15, CAO16, CAO17, CAO18, CAO19, CAO20, CAO21, CAO22, CAO23, CAO24
, CBI1, CBI2, CBI3, CBI4, CBI5, CBI6, CBI7, CBI8, CBI9, CBI10, CBI11, CBI12, CBI13, CBI14, CBI15, CBI16, CBI17, CBI18, CBO1, CBO2, CBO3
, CBO4, CBO5, CBO6, CBO7, CBO8, CBO9, CBO10, CBO11, CBO12, CBO13, CBO14, CBO15, CBO16, CBO17, CBO18, CCI, CCO, CI, CK, CO43, CO57
, RESERVED, CZI1, CZI2, CZI3, CZI4, CZI5, CZI6, CZI7, CZI8, CZI9, CZI10, CZI11, CZI12, CZI13, CZI14, CZI15, CZI16, CZI17, CZI18, CZI19, CZI20
, CZI21, CZI22, CZI23, CZI24, CZI25, CZI26, CZI27, CZI28, CZI29, CZI30, CZI31, CZI32, CZI33, CZI34, CZI35, CZI36, CZI37, CZI38, CZI39, CZI40, CZI41
, CZI42, CZI43, CZI44, CZI45, CZI46, CZI47, CZI48, CZI49, CZI50, CZI51, CZI52, CZI53, CZI54, CZI55, CZI56, CZO1, CZO2, CZO3, CZO4, CZO5, CZO6
, CZO7, CZO8, CZO9, CZO10, CZO11, CZO12, CZO13, CZO14, CZO15, CZO16, CZO17, CZO18, CZO19, CZO20, CZO21, CZO22, CZO23, CZO24, CZO25, CZO26, CZO27
, CZO28, CZO29, CZO30, CZO31, CZO32, CZO33, CZO34, CZO35, CZO36, CZO37, CZO38, CZO39, CZO40, CZO41, CZO42, CZO43, CZO44, CZO45, CZO46, CZO47, CZO48
, CZO49, CZO50, CZO51, CZO52, CZO53, CZO54, CZO55, CZO56, D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13
, D14, D15, D16, D17, D18, OVF, R, RZ, WE, WEZ, Z1, Z2, Z3, Z4, Z5, Z6, Z7, Z8, Z9, Z10, Z11
, Z12, Z13, Z14, Z15, Z16, Z17, Z18, Z19, Z20, Z21, Z22, Z23, Z24, Z25, Z26, Z27, Z28, Z29, Z30, Z31, Z32
, Z33, Z34, Z35, Z36, Z37, Z38, Z39, Z40, Z41, Z42, Z43, Z44, Z45, Z46, Z47, Z48, Z49, Z50, Z51, Z52, Z53
, Z54, Z55, Z56);
    input A1;
    input A10;
    input A11;
    input A12;
    input A13;
    input A14;
    input A15;
    input A16;
    input A17;
    input A18;
    input A19;
    input A2;
    input A20;
    input A21;
    input A22;
    input A23;
    input A24;
    input A3;
    input A4;
    input A5;
    input A6;
    input A7;
    input A8;
    input A9;
    input B1;
    input B10;
    input B11;
    input B12;
    input B13;
    input B14;
    input B15;
    input B16;
    input B17;
    input B18;
    input B2;
    input B3;
    input B4;
    input B5;
    input B6;
    input B7;
    input B8;
    input B9;
    input C1;
    input C10;
    input C11;
    input C12;
    input C13;
    input C14;
    input C15;
    input C16;
    input C17;
    input C18;
    input C19;
    input C2;
    input C20;
    input C21;
    input C22;
    input C23;
    input C24;
    input C25;
    input C26;
    input C27;
    input C28;
    input C29;
    input C3;
    input C30;
    input C31;
    input C32;
    input C33;
    input C34;
    input C35;
    input C36;
    input C4;
    input C5;
    input C6;
    input C7;
    input C8;
    input C9;
    input CAI1;
    input CAI10;
    input CAI11;
    input CAI12;
    input CAI13;
    input CAI14;
    input CAI15;
    input CAI16;
    input CAI17;
    input CAI18;
    input CAI19;
    input CAI2;
    input CAI20;
    input CAI21;
    input CAI22;
    input CAI23;
    input CAI24;
    input CAI3;
    input CAI4;
    input CAI5;
    input CAI6;
    input CAI7;
    input CAI8;
    input CAI9;
    output CAO1;
    output CAO10;
    output CAO11;
    output CAO12;
    output CAO13;
    output CAO14;
    output CAO15;
    output CAO16;
    output CAO17;
    output CAO18;
    output CAO19;
    output CAO2;
    output CAO20;
    output CAO21;
    output CAO22;
    output CAO23;
    output CAO24;
    output CAO3;
    output CAO4;
    output CAO5;
    output CAO6;
    output CAO7;
    output CAO8;
    output CAO9;
    input CBI1;
    input CBI10;
    input CBI11;
    input CBI12;
    input CBI13;
    input CBI14;
    input CBI15;
    input CBI16;
    input CBI17;
    input CBI18;
    input CBI2;
    input CBI3;
    input CBI4;
    input CBI5;
    input CBI6;
    input CBI7;
    input CBI8;
    input CBI9;
    output CBO1;
    output CBO10;
    output CBO11;
    output CBO12;
    output CBO13;
    output CBO14;
    output CBO15;
    output CBO16;
    output CBO17;
    output CBO18;
    output CBO2;
    output CBO3;
    output CBO4;
    output CBO5;
    output CBO6;
    output CBO7;
    output CBO8;
    output CBO9;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO43;
    output CO57;
    input CZI1;
    input CZI10;
    input CZI11;
    input CZI12;
    input CZI13;
    input CZI14;
    input CZI15;
    input CZI16;
    input CZI17;
    input CZI18;
    input CZI19;
    input CZI2;
    input CZI20;
    input CZI21;
    input CZI22;
    input CZI23;
    input CZI24;
    input CZI25;
    input CZI26;
    input CZI27;
    input CZI28;
    input CZI29;
    input CZI3;
    input CZI30;
    input CZI31;
    input CZI32;
    input CZI33;
    input CZI34;
    input CZI35;
    input CZI36;
    input CZI37;
    input CZI38;
    input CZI39;
    input CZI4;
    input CZI40;
    input CZI41;
    input CZI42;
    input CZI43;
    input CZI44;
    input CZI45;
    input CZI46;
    input CZI47;
    input CZI48;
    input CZI49;
    input CZI5;
    input CZI50;
    input CZI51;
    input CZI52;
    input CZI53;
    input CZI54;
    input CZI55;
    input CZI56;
    input CZI6;
    input CZI7;
    input CZI8;
    input CZI9;
    output CZO1;
    output CZO10;
    output CZO11;
    output CZO12;
    output CZO13;
    output CZO14;
    output CZO15;
    output CZO16;
    output CZO17;
    output CZO18;
    output CZO19;
    output CZO2;
    output CZO20;
    output CZO21;
    output CZO22;
    output CZO23;
    output CZO24;
    output CZO25;
    output CZO26;
    output CZO27;
    output CZO28;
    output CZO29;
    output CZO3;
    output CZO30;
    output CZO31;
    output CZO32;
    output CZO33;
    output CZO34;
    output CZO35;
    output CZO36;
    output CZO37;
    output CZO38;
    output CZO39;
    output CZO4;
    output CZO40;
    output CZO41;
    output CZO42;
    output CZO43;
    output CZO44;
    output CZO45;
    output CZO46;
    output CZO47;
    output CZO48;
    output CZO49;
    output CZO5;
    output CZO50;
    output CZO51;
    output CZO52;
    output CZO53;
    output CZO54;
    output CZO55;
    output CZO56;
    output CZO6;
    output CZO7;
    output CZO8;
    output CZO9;
    input D1;
    input D10;
    input D11;
    input D12;
    input D13;
    input D14;
    input D15;
    input D16;
    input D17;
    input D18;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input D7;
    input D8;
    input D9;
    output OVF;
    input R;
    output RESERVED;
    input RZ;
    input WE;
    input WEZ;
    output Z1;
    output Z10;
    output Z11;
    output Z12;
    output Z13;
    output Z14;
    output Z15;
    output Z16;
    output Z17;
    output Z18;
    output Z19;
    output Z2;
    output Z20;
    output Z21;
    output Z22;
    output Z23;
    output Z24;
    output Z25;
    output Z26;
    output Z27;
    output Z28;
    output Z29;
    output Z3;
    output Z30;
    output Z31;
    output Z32;
    output Z33;
    output Z34;
    output Z35;
    output Z36;
    output Z37;
    output Z38;
    output Z39;
    output Z4;
    output Z40;
    output Z41;
    output Z42;
    output Z43;
    output Z44;
    output Z45;
    output Z46;
    output Z47;
    output Z48;
    output Z49;
    output Z5;
    output Z50;
    output Z51;
    output Z52;
    output Z53;
    output Z54;
    output Z55;
    output Z56;
    output Z6;
    output Z7;
    output Z8;
    output Z9;
    parameter raw_config0 = 27'b000000000000000000000000000;
    parameter raw_config1 = 24'b000000000000000000000000;
    parameter raw_config2 = 14'b00000000000000;
    parameter raw_config3 = 3'b000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_DSP_U_SPLIT(CK, R, RZ, WE, WEZ, CI, CCI, CO42, CO56, OVF, CCO, A, B, C, D, Z, CAI, CBI, CZI, CAO, CBO
, CZO);
    input [23:0] A;
    input [17:0] B;
    input [35:0] C;
    input [23:0] CAI;
    output [23:0] CAO;
    input [17:0] CBI;
    output [17:0] CBO;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO42;
    output CO56;
    input [55:0] CZI;
    output [55:0] CZO;
    input [17:0] D;
    output OVF;
    input R;
    input RZ;
    input WE;
    input WEZ;
    output [55:0] Z;
    parameter ALU_DYNAMIC_OP = 2'b00;
    parameter ALU_OP = 3'b000;
    parameter ENABLE_PR_A_RST = 1'b0;
    parameter ENABLE_PR_B_RST = 1'b0;
    parameter ENABLE_PR_CCO_RST = 1'b0;
    parameter ENABLE_PR_CI_RST = 1'b0;
    parameter ENABLE_PR_CO_RST = 1'b0;
    parameter ENABLE_PR_CZ_RST = 1'b0;
    parameter ENABLE_PR_C_RST = 1'b0;
    parameter ENABLE_PR_D_RST = 1'b0;
    parameter ENABLE_PR_MULT_RST = 1'b0;
    parameter ENABLE_PR_OV_RST = 1'b0;
    parameter ENABLE_PR_P_RST = 1'b0;
    parameter ENABLE_PR_X_RST = 1'b0;
    parameter ENABLE_PR_Y_RST = 1'b0;
    parameter ENABLE_PR_Z_RST = 1'b0;
    parameter ENABLE_SATURATION = 1'b0;
    parameter INV_RST = 1'b0;
    parameter INV_RSTZ = 1'b0;
    parameter INV_WE = 1'b0;
    parameter INV_WEZ = 1'b0;
    parameter MUX_A = 1'b0;
    parameter MUX_B = 1'b0;
    parameter MUX_CCI = 1'b0;
    parameter MUX_CCO = 1'b0;
    parameter MUX_CI = 1'b0;
    parameter MUX_CZ = 1'b0;
    parameter MUX_P = 1'b0;
    parameter MUX_X = 3'b000;
    parameter MUX_Y = 1'b0;
    parameter MUX_Z = 1'b0;
    parameter PRE_ADDER_OP = 1'b0;
    parameter PR_A_CASCADE_MUX = 2'b00;
    parameter PR_A_MUX = 2'b00;
    parameter PR_B_CASCADE_MUX = 2'b00;
    parameter PR_B_MUX = 2'b00;
    parameter PR_CCO_MUX = 1'b0;
    parameter PR_CI_MUX = 1'b0;
    parameter PR_CO_MUX = 1'b0;
    parameter PR_CZ_MUX = 1'b0;
    parameter PR_C_MUX = 1'b0;
    parameter PR_D_MUX = 1'b0;
    parameter PR_MULT_MUX = 1'b0;
    parameter PR_OV_MUX = 1'b0;
    parameter PR_P_MUX = 1'b0;
    parameter PR_RSTZ_MUX = 1'b0;
    parameter PR_RST_MUX = 1'b0;
    parameter PR_WEZ_MUX = 1'b0;
    parameter PR_WE_MUX = 1'b0;
    parameter PR_X_MUX = 1'b0;
    parameter PR_Y_MUX = 1'b0;
    parameter PR_Z_MUX = 1'b0;
    parameter SATURATION_RANK = 6'b000000;
    parameter SIGNED_MODE = 1'b0;
endmodule

(* blackbox *)
module NX_DSP_U_WRAP(CCI, CCO, CI, CK, CO43, CO57, OVF, R, RZ, WE, WEZ, A, B, C, D, Z, CAI, CBI, CZI, CAO, CBO
, CZO);
    input [23:0] A;
    input [17:0] B;
    input [35:0] C;
    input [23:0] CAI;
    output [23:0] CAO;
    input [17:0] CBI;
    output [17:0] CBO;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO43;
    output CO57;
    input [55:0] CZI;
    output [55:0] CZO;
    input [17:0] D;
    output OVF;
    input R;
    input RZ;
    input WE;
    input WEZ;
    output [55:0] Z;
    parameter raw_config0 = 27'b000000000000000000000000000;
    parameter raw_config1 = 24'b000000000000000000000000;
    parameter raw_config2 = 14'b00000000000000;
    parameter raw_config3 = 3'b000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_DSP_WRAP(CCI, CCO, CI, CK, CO, CO37, CO49, OVF, R, RZ, WE, A, B, C, D, Z, CAI, CBI, CZI, CAO, CBO
, CZO);
    input [23:0] A;
    input [17:0] B;
    input [35:0] C;
    input [17:0] CAI;
    output [17:0] CAO;
    input [17:0] CBI;
    output [17:0] CBO;
    input CCI;
    output CCO;
    input CI;
    input CK;
    output CO;
    output CO37;
    output CO49;
    input [55:0] CZI;
    output [55:0] CZO;
    input [17:0] D;
    output OVF;
    input R;
    input RZ;
    input WE;
    output [55:0] Z;
    parameter raw_config0 = 20'b00000000000000000000;
    parameter raw_config1 = 19'b0000000000000000000;
    parameter raw_config2 = 13'b0000000000000;
    parameter raw_config3 = 7'b0000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_ECC(CKD, CHK, COR, ERR);
    input CHK;
    input CKD;
    output COR;
    output ERR;
endmodule

(* blackbox *)
module NX_FIFO_DPREG(RCK, WCK, WE, WEA, WRSTI, WRSTO, WEQ, RRSTI, RRSTO, REQ, I, O, WAI, WAO, RAI, RAO);
    input [17:0] I;
    output [17:0] O;
    input [5:0] RAI;
    output [5:0] RAO;
    input RCK;
    output REQ;
    input RRSTI;
    output RRSTO;
    input [5:0] WAI;
    output [5:0] WAO;
    input WCK;
    input WE;
    input WEA;
    output WEQ;
    input WRSTI;
    output WRSTO;
    parameter rck_edge = 1'b0;
    parameter read_addr_inv = 6'b000000;
    parameter use_read_arst = 1'b0;
    parameter use_write_arst = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_FIFO_U(RCK, WCK, WE, WEA, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17
, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, I32, I33, I34, I35, I36, O1, O2
, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23
, O24, O25, O26, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, WRSTI, WAI1, WAI2, WAI3, WAI4, WAI5, WAI6, WAI7
, WRSTO, WAO1, WAO2, WAO3, WAO4, WAO5, WAO6, WAO7, WEQ1, WEQ2, RRSTI, RAI1, RAI2, RAI3, RAI4, RAI5, RAI6, RAI7, RRSTO, RAO1, RAO2
, RAO3, RAO4, RAO5, RAO6, RAO7, REQ1, REQ2);
    input I1;
    input I10;
    input I11;
    input I12;
    input I13;
    input I14;
    input I15;
    input I16;
    input I17;
    input I18;
    input I19;
    input I2;
    input I20;
    input I21;
    input I22;
    input I23;
    input I24;
    input I25;
    input I26;
    input I27;
    input I28;
    input I29;
    input I3;
    input I30;
    input I31;
    input I32;
    input I33;
    input I34;
    input I35;
    input I36;
    input I4;
    input I5;
    input I6;
    input I7;
    input I8;
    input I9;
    output O1;
    output O10;
    output O11;
    output O12;
    output O13;
    output O14;
    output O15;
    output O16;
    output O17;
    output O18;
    output O19;
    output O2;
    output O20;
    output O21;
    output O22;
    output O23;
    output O24;
    output O25;
    output O26;
    output O27;
    output O28;
    output O29;
    output O3;
    output O30;
    output O31;
    output O32;
    output O33;
    output O34;
    output O35;
    output O36;
    output O4;
    output O5;
    output O6;
    output O7;
    output O8;
    output O9;
    input RAI1;
    input RAI2;
    input RAI3;
    input RAI4;
    input RAI5;
    input RAI6;
    input RAI7;
    output RAO1;
    output RAO2;
    output RAO3;
    output RAO4;
    output RAO5;
    output RAO6;
    output RAO7;
    input RCK;
    output REQ1;
    output REQ2;
    input RRSTI;
    output RRSTO;
    input WAI1;
    input WAI2;
    input WAI3;
    input WAI4;
    input WAI5;
    input WAI6;
    input WAI7;
    output WAO1;
    output WAO2;
    output WAO3;
    output WAO4;
    output WAO5;
    output WAO6;
    output WAO7;
    input WCK;
    input WE;
    input WEA;
    output WEQ1;
    output WEQ2;
    input WRSTI;
    output WRSTO;
    parameter mode = 0;
    parameter rck_edge = 1'b0;
    parameter read_addr_inv = 7'b0000000;
    parameter use_read_arst = 1'b0;
    parameter use_write_arst = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_HSSL_L_FULL(hssl_clk_user_i, hssl_clk_ref_i, hssl_clock_o, usr_com_tx_pma_pre_sign_i, usr_com_tx_pma_pre_en_i, usr_com_tx_pma_main_sign_i, usr_com_rx_pma_m_eye_i, usr_com_tx_pma_post_sign_i, usr_pll_pma_rst_n_i, usr_main_rst_n_i, usr_calibrate_pma_en_i, usr_pcs_ctrl_pll_lock_en_i, usr_pcs_ctrl_ovs_en_i, usr_pll_lock_o, usr_calibrate_pma_out_o, pma_clk_ext_i, usr_tx0_ctrl_replace_en_i, usr_tx0_rst_n_i, usr_tx0_pma_clk_en_i, usr_tx0_busy_o, pma_tx0_o
, usr_rx0_ctrl_dscr_en_i, usr_rx0_ctrl_dec_en_i, usr_rx0_ctrl_align_en_i, usr_rx0_ctrl_align_sync_i, usr_rx0_ctrl_replace_en_i, usr_rx0_ctrl_el_buff_rst_i, usr_rx0_ctrl_el_buff_fifo_en_i, usr_rx0_rst_n_i, usr_rx0_pma_cdr_rst_i, usr_rx0_pma_ckgen_rst_n_i, usr_rx0_pma_pll_rst_n_i, usr_rx0_pma_loss_of_signal_o, usr_rx0_ctrl_char_is_aligned_o, usr_rx0_busy_o, usr_rx0_pll_lock_o, pma_rx0_i, usr_tx1_ctrl_replace_en_i, usr_tx1_rst_n_i, usr_tx1_pma_clk_en_i, usr_tx1_busy_o, pma_tx1_o
, usr_rx1_ctrl_dscr_en_i, usr_rx1_ctrl_dec_en_i, usr_rx1_ctrl_align_en_i, usr_rx1_ctrl_align_sync_i, usr_rx1_ctrl_replace_en_i, usr_rx1_ctrl_el_buff_rst_i, usr_rx1_ctrl_el_buff_fifo_en_i, usr_rx1_rst_n_i, usr_rx1_pma_cdr_rst_i, usr_rx1_pma_ckgen_rst_n_i, usr_rx1_pma_pll_rst_n_i, usr_rx1_pma_loss_of_signal_o, usr_rx1_ctrl_char_is_aligned_o, usr_rx1_busy_o, usr_rx1_pll_lock_o, pma_rx1_i, usr_tx2_ctrl_replace_en_i, usr_tx2_rst_n_i, usr_tx2_pma_clk_en_i, usr_tx2_busy_o, pma_tx2_o
, usr_rx2_ctrl_dscr_en_i, usr_rx2_ctrl_dec_en_i, usr_rx2_ctrl_align_en_i, usr_rx2_ctrl_align_sync_i, usr_rx2_ctrl_replace_en_i, usr_rx2_ctrl_el_buff_rst_i, usr_rx2_ctrl_el_buff_fifo_en_i, usr_rx2_rst_n_i, usr_rx2_pma_cdr_rst_i, usr_rx2_pma_ckgen_rst_n_i, usr_rx2_pma_pll_rst_n_i, usr_rx2_pma_loss_of_signal_o, usr_rx2_ctrl_char_is_aligned_o, usr_rx2_busy_o, usr_rx2_pll_lock_o, pma_rx2_i, usr_tx3_ctrl_replace_en_i, usr_tx3_rst_n_i, usr_tx3_pma_clk_en_i, usr_tx3_busy_o, pma_tx3_o
, usr_rx3_ctrl_dscr_en_i, usr_rx3_ctrl_dec_en_i, usr_rx3_ctrl_align_en_i, usr_rx3_ctrl_align_sync_i, usr_rx3_ctrl_replace_en_i, usr_rx3_ctrl_el_buff_rst_i, usr_rx3_ctrl_el_buff_fifo_en_i, usr_rx3_rst_n_i, usr_rx3_pma_cdr_rst_i, usr_rx3_pma_ckgen_rst_n_i, usr_rx3_pma_pll_rst_n_i, usr_rx3_pma_loss_of_signal_o, usr_rx3_ctrl_char_is_aligned_o, usr_rx3_busy_o, usr_rx3_pll_lock_o, pma_rx3_i, usr_tx4_ctrl_replace_en_i, usr_tx4_rst_n_i, usr_tx4_pma_clk_en_i, usr_tx4_busy_o, pma_tx4_o
, usr_rx4_ctrl_dscr_en_i, usr_rx4_ctrl_dec_en_i, usr_rx4_ctrl_align_en_i, usr_rx4_ctrl_align_sync_i, usr_rx4_ctrl_replace_en_i, usr_rx4_ctrl_el_buff_rst_i, usr_rx4_ctrl_el_buff_fifo_en_i, usr_rx4_rst_n_i, usr_rx4_pma_cdr_rst_i, usr_rx4_pma_ckgen_rst_n_i, usr_rx4_pma_pll_rst_n_i, usr_rx4_pma_loss_of_signal_o, usr_rx4_ctrl_char_is_aligned_o, usr_rx4_busy_o, usr_rx4_pll_lock_o, pma_rx4_i, usr_tx5_ctrl_replace_en_i, usr_tx5_rst_n_i, usr_tx5_pma_clk_en_i, usr_tx5_busy_o, pma_tx5_o
, usr_rx5_ctrl_dscr_en_i, usr_rx5_ctrl_dec_en_i, usr_rx5_ctrl_align_en_i, usr_rx5_ctrl_align_sync_i, usr_rx5_ctrl_replace_en_i, usr_rx5_ctrl_el_buff_rst_i, usr_rx5_ctrl_el_buff_fifo_en_i, usr_rx5_rst_n_i, usr_rx5_pma_cdr_rst_i, usr_rx5_pma_ckgen_rst_n_i, usr_rx5_pma_pll_rst_n_i, usr_rx5_pma_loss_of_signal_o, usr_rx5_ctrl_char_is_aligned_o, usr_rx5_busy_o, usr_rx5_pll_lock_o, pma_rx5_i, usr_com_tx_pma_main_en_i, usr_com_tx_pma_margin_sel_i, usr_com_tx_pma_margin_input_sel_i, usr_com_tx_pma_margin_sel_var_i, usr_com_tx_pma_margin_input_sel_var_i
, usr_com_tx_pma_post_en_i, usr_com_tx_pma_post_input_sel_i, usr_com_tx_pma_post_input_sel_var_i, usr_com_rx_pma_ctle_cap_i, usr_com_rx_pma_ctle_resp_i, usr_com_rx_pma_ctle_resn_i, usr_com_ctrl_tx_sel_i, usr_com_ctrl_rx_sel_i, usr_calibrate_pma_res_p1_i, usr_calibrate_pma_res_n2_i, usr_calibrate_pma_res_n3_i, usr_calibrate_pma_res_p4_i, usr_calibrate_pma_sel_i, usr_main_test_i, usr_main_test_o, usr_tx0_ctrl_enc_en_i, usr_tx0_ctrl_char_is_k_i, usr_tx0_ctrl_scr_en_i, usr_tx0_ctrl_end_of_multiframe_i, usr_tx0_ctrl_end_of_frame_i, usr_tx0_test_i
, usr_tx0_data_i, usr_tx0_test_o, usr_rx0_data_o, usr_rx0_ctrl_ovs_bit_sel_i, usr_rx0_test_i, usr_rx0_ctrl_char_is_comma_o, usr_rx0_ctrl_char_is_k_o, usr_rx0_ctrl_not_in_table_o, usr_rx0_ctrl_disp_err_o, usr_rx0_ctrl_char_is_a_o, usr_rx0_ctrl_char_is_f_o, usr_rx0_test_o, usr_tx1_ctrl_enc_en_i, usr_tx1_ctrl_char_is_k_i, usr_tx1_ctrl_scr_en_i, usr_tx1_ctrl_end_of_multiframe_i, usr_tx1_ctrl_end_of_frame_i, usr_tx1_test_i, usr_tx1_data_i, usr_tx1_test_o, usr_rx1_data_o
, usr_rx1_ctrl_ovs_bit_sel_i, usr_rx1_test_i, usr_rx1_ctrl_char_is_comma_o, usr_rx1_ctrl_char_is_k_o, usr_rx1_ctrl_not_in_table_o, usr_rx1_ctrl_disp_err_o, usr_rx1_ctrl_char_is_a_o, usr_rx1_ctrl_char_is_f_o, usr_rx1_test_o, usr_tx2_ctrl_enc_en_i, usr_tx2_ctrl_char_is_k_i, usr_tx2_ctrl_scr_en_i, usr_tx2_ctrl_end_of_multiframe_i, usr_tx2_ctrl_end_of_frame_i, usr_tx2_test_i, usr_tx2_data_i, usr_tx2_test_o, usr_rx2_data_o, usr_rx2_ctrl_ovs_bit_sel_i, usr_rx2_test_i, usr_rx2_ctrl_char_is_comma_o
, usr_rx2_ctrl_char_is_k_o, usr_rx2_ctrl_not_in_table_o, usr_rx2_ctrl_disp_err_o, usr_rx2_ctrl_char_is_a_o, usr_rx2_ctrl_char_is_f_o, usr_rx2_test_o, usr_tx3_ctrl_enc_en_i, usr_tx3_ctrl_char_is_k_i, usr_tx3_ctrl_scr_en_i, usr_tx3_ctrl_end_of_multiframe_i, usr_tx3_ctrl_end_of_frame_i, usr_tx3_test_i, usr_tx3_data_i, usr_tx3_test_o, usr_rx3_data_o, usr_rx3_ctrl_ovs_bit_sel_i, usr_rx3_test_i, usr_rx3_ctrl_char_is_comma_o, usr_rx3_ctrl_char_is_k_o, usr_rx3_ctrl_not_in_table_o, usr_rx3_ctrl_disp_err_o
, usr_rx3_ctrl_char_is_a_o, usr_rx3_ctrl_char_is_f_o, usr_rx3_test_o, usr_tx4_ctrl_enc_en_i, usr_tx4_ctrl_char_is_k_i, usr_tx4_ctrl_scr_en_i, usr_tx4_ctrl_end_of_multiframe_i, usr_tx4_ctrl_end_of_frame_i, usr_tx4_test_i, usr_tx4_data_i, usr_tx4_test_o, usr_rx4_data_o, usr_rx4_ctrl_ovs_bit_sel_i, usr_rx4_test_i, usr_rx4_ctrl_char_is_comma_o, usr_rx4_ctrl_char_is_k_o, usr_rx4_ctrl_not_in_table_o, usr_rx4_ctrl_disp_err_o, usr_rx4_ctrl_char_is_a_o, usr_rx4_ctrl_char_is_f_o, usr_rx4_test_o
, usr_tx5_ctrl_enc_en_i, usr_tx5_ctrl_char_is_k_i, usr_tx5_ctrl_scr_en_i, usr_tx5_ctrl_end_of_multiframe_i, usr_tx5_ctrl_end_of_frame_i, usr_tx5_test_i, usr_tx5_data_i, usr_tx5_test_o, usr_rx5_data_o, usr_rx5_ctrl_ovs_bit_sel_i, usr_rx5_test_i, usr_rx5_ctrl_char_is_comma_o, usr_rx5_ctrl_char_is_k_o, usr_rx5_ctrl_not_in_table_o, usr_rx5_ctrl_disp_err_o, usr_rx5_ctrl_char_is_a_o, usr_rx5_ctrl_char_is_f_o, usr_rx5_test_o, usr_com_tx_pma_pre_input_sel_i);
    input hssl_clk_ref_i;
    input hssl_clk_user_i;
    output hssl_clock_o;
    input pma_clk_ext_i;
    input pma_rx0_i;
    input pma_rx1_i;
    input pma_rx2_i;
    input pma_rx3_i;
    input pma_rx4_i;
    input pma_rx5_i;
    output pma_tx0_o;
    output pma_tx1_o;
    output pma_tx2_o;
    output pma_tx3_o;
    output pma_tx4_o;
    output pma_tx5_o;
    input usr_calibrate_pma_en_i;
    output usr_calibrate_pma_out_o;
    input [7:0] usr_calibrate_pma_res_n2_i;
    input [7:0] usr_calibrate_pma_res_n3_i;
    input [7:0] usr_calibrate_pma_res_p1_i;
    input [7:0] usr_calibrate_pma_res_p4_i;
    input [3:0] usr_calibrate_pma_sel_i;
    input [5:0] usr_com_ctrl_rx_sel_i;
    input [5:0] usr_com_ctrl_tx_sel_i;
    input [3:0] usr_com_rx_pma_ctle_cap_i;
    input [3:0] usr_com_rx_pma_ctle_resn_i;
    input [3:0] usr_com_rx_pma_ctle_resp_i;
    input usr_com_rx_pma_m_eye_i;
    input [5:0] usr_com_tx_pma_main_en_i;
    input usr_com_tx_pma_main_sign_i;
    input [3:0] usr_com_tx_pma_margin_input_sel_i;
    input [4:0] usr_com_tx_pma_margin_input_sel_var_i;
    input [3:0] usr_com_tx_pma_margin_sel_i;
    input [4:0] usr_com_tx_pma_margin_sel_var_i;
    input [4:0] usr_com_tx_pma_post_en_i;
    input [3:0] usr_com_tx_pma_post_input_sel_i;
    input [3:0] usr_com_tx_pma_post_input_sel_var_i;
    input usr_com_tx_pma_post_sign_i;
    input usr_com_tx_pma_pre_en_i;
    input [3:0] usr_com_tx_pma_pre_input_sel_i;
    input usr_com_tx_pma_pre_sign_i;
    input usr_main_rst_n_i;
    input [7:0] usr_main_test_i;
    output [7:0] usr_main_test_o;
    input usr_pcs_ctrl_ovs_en_i;
    input usr_pcs_ctrl_pll_lock_en_i;
    output usr_pll_lock_o;
    input usr_pll_pma_rst_n_i;
    output usr_rx0_busy_o;
    input usr_rx0_ctrl_align_en_i;
    input usr_rx0_ctrl_align_sync_i;
    output [7:0] usr_rx0_ctrl_char_is_a_o;
    output usr_rx0_ctrl_char_is_aligned_o;
    output [7:0] usr_rx0_ctrl_char_is_comma_o;
    output [7:0] usr_rx0_ctrl_char_is_f_o;
    output [7:0] usr_rx0_ctrl_char_is_k_o;
    input usr_rx0_ctrl_dec_en_i;
    output [7:0] usr_rx0_ctrl_disp_err_o;
    input usr_rx0_ctrl_dscr_en_i;
    input usr_rx0_ctrl_el_buff_fifo_en_i;
    input usr_rx0_ctrl_el_buff_rst_i;
    output [7:0] usr_rx0_ctrl_not_in_table_o;
    input [1:0] usr_rx0_ctrl_ovs_bit_sel_i;
    input usr_rx0_ctrl_replace_en_i;
    output [63:0] usr_rx0_data_o;
    output usr_rx0_pll_lock_o;
    input usr_rx0_pma_cdr_rst_i;
    input usr_rx0_pma_ckgen_rst_n_i;
    output usr_rx0_pma_loss_of_signal_o;
    input usr_rx0_pma_pll_rst_n_i;
    input usr_rx0_rst_n_i;
    input [3:0] usr_rx0_test_i;
    output [7:0] usr_rx0_test_o;
    output usr_rx1_busy_o;
    input usr_rx1_ctrl_align_en_i;
    input usr_rx1_ctrl_align_sync_i;
    output [7:0] usr_rx1_ctrl_char_is_a_o;
    output usr_rx1_ctrl_char_is_aligned_o;
    output [7:0] usr_rx1_ctrl_char_is_comma_o;
    output [7:0] usr_rx1_ctrl_char_is_f_o;
    output [7:0] usr_rx1_ctrl_char_is_k_o;
    input usr_rx1_ctrl_dec_en_i;
    output [7:0] usr_rx1_ctrl_disp_err_o;
    input usr_rx1_ctrl_dscr_en_i;
    input usr_rx1_ctrl_el_buff_fifo_en_i;
    input usr_rx1_ctrl_el_buff_rst_i;
    output [7:0] usr_rx1_ctrl_not_in_table_o;
    input [1:0] usr_rx1_ctrl_ovs_bit_sel_i;
    input usr_rx1_ctrl_replace_en_i;
    output [63:0] usr_rx1_data_o;
    output usr_rx1_pll_lock_o;
    input usr_rx1_pma_cdr_rst_i;
    input usr_rx1_pma_ckgen_rst_n_i;
    output usr_rx1_pma_loss_of_signal_o;
    input usr_rx1_pma_pll_rst_n_i;
    input usr_rx1_rst_n_i;
    input [3:0] usr_rx1_test_i;
    output [7:0] usr_rx1_test_o;
    output usr_rx2_busy_o;
    input usr_rx2_ctrl_align_en_i;
    input usr_rx2_ctrl_align_sync_i;
    output [7:0] usr_rx2_ctrl_char_is_a_o;
    output usr_rx2_ctrl_char_is_aligned_o;
    output [7:0] usr_rx2_ctrl_char_is_comma_o;
    output [7:0] usr_rx2_ctrl_char_is_f_o;
    output [7:0] usr_rx2_ctrl_char_is_k_o;
    input usr_rx2_ctrl_dec_en_i;
    output [7:0] usr_rx2_ctrl_disp_err_o;
    input usr_rx2_ctrl_dscr_en_i;
    input usr_rx2_ctrl_el_buff_fifo_en_i;
    input usr_rx2_ctrl_el_buff_rst_i;
    output [7:0] usr_rx2_ctrl_not_in_table_o;
    input [1:0] usr_rx2_ctrl_ovs_bit_sel_i;
    input usr_rx2_ctrl_replace_en_i;
    output [63:0] usr_rx2_data_o;
    output usr_rx2_pll_lock_o;
    input usr_rx2_pma_cdr_rst_i;
    input usr_rx2_pma_ckgen_rst_n_i;
    output usr_rx2_pma_loss_of_signal_o;
    input usr_rx2_pma_pll_rst_n_i;
    input usr_rx2_rst_n_i;
    input [3:0] usr_rx2_test_i;
    output [7:0] usr_rx2_test_o;
    output usr_rx3_busy_o;
    input usr_rx3_ctrl_align_en_i;
    input usr_rx3_ctrl_align_sync_i;
    output [7:0] usr_rx3_ctrl_char_is_a_o;
    output usr_rx3_ctrl_char_is_aligned_o;
    output [7:0] usr_rx3_ctrl_char_is_comma_o;
    output [7:0] usr_rx3_ctrl_char_is_f_o;
    output [7:0] usr_rx3_ctrl_char_is_k_o;
    input usr_rx3_ctrl_dec_en_i;
    output [7:0] usr_rx3_ctrl_disp_err_o;
    input usr_rx3_ctrl_dscr_en_i;
    input usr_rx3_ctrl_el_buff_fifo_en_i;
    input usr_rx3_ctrl_el_buff_rst_i;
    output [7:0] usr_rx3_ctrl_not_in_table_o;
    input [1:0] usr_rx3_ctrl_ovs_bit_sel_i;
    input usr_rx3_ctrl_replace_en_i;
    output [63:0] usr_rx3_data_o;
    output usr_rx3_pll_lock_o;
    input usr_rx3_pma_cdr_rst_i;
    input usr_rx3_pma_ckgen_rst_n_i;
    output usr_rx3_pma_loss_of_signal_o;
    input usr_rx3_pma_pll_rst_n_i;
    input usr_rx3_rst_n_i;
    input [3:0] usr_rx3_test_i;
    output [7:0] usr_rx3_test_o;
    output usr_rx4_busy_o;
    input usr_rx4_ctrl_align_en_i;
    input usr_rx4_ctrl_align_sync_i;
    output [7:0] usr_rx4_ctrl_char_is_a_o;
    output usr_rx4_ctrl_char_is_aligned_o;
    output [7:0] usr_rx4_ctrl_char_is_comma_o;
    output [7:0] usr_rx4_ctrl_char_is_f_o;
    output [7:0] usr_rx4_ctrl_char_is_k_o;
    input usr_rx4_ctrl_dec_en_i;
    output [7:0] usr_rx4_ctrl_disp_err_o;
    input usr_rx4_ctrl_dscr_en_i;
    input usr_rx4_ctrl_el_buff_fifo_en_i;
    input usr_rx4_ctrl_el_buff_rst_i;
    output [7:0] usr_rx4_ctrl_not_in_table_o;
    input [1:0] usr_rx4_ctrl_ovs_bit_sel_i;
    input usr_rx4_ctrl_replace_en_i;
    output [63:0] usr_rx4_data_o;
    output usr_rx4_pll_lock_o;
    input usr_rx4_pma_cdr_rst_i;
    input usr_rx4_pma_ckgen_rst_n_i;
    output usr_rx4_pma_loss_of_signal_o;
    input usr_rx4_pma_pll_rst_n_i;
    input usr_rx4_rst_n_i;
    input [3:0] usr_rx4_test_i;
    output [7:0] usr_rx4_test_o;
    output usr_rx5_busy_o;
    input usr_rx5_ctrl_align_en_i;
    input usr_rx5_ctrl_align_sync_i;
    output [7:0] usr_rx5_ctrl_char_is_a_o;
    output usr_rx5_ctrl_char_is_aligned_o;
    output [7:0] usr_rx5_ctrl_char_is_comma_o;
    output [7:0] usr_rx5_ctrl_char_is_f_o;
    output [7:0] usr_rx5_ctrl_char_is_k_o;
    input usr_rx5_ctrl_dec_en_i;
    output [7:0] usr_rx5_ctrl_disp_err_o;
    input usr_rx5_ctrl_dscr_en_i;
    input usr_rx5_ctrl_el_buff_fifo_en_i;
    input usr_rx5_ctrl_el_buff_rst_i;
    output [7:0] usr_rx5_ctrl_not_in_table_o;
    input [1:0] usr_rx5_ctrl_ovs_bit_sel_i;
    input usr_rx5_ctrl_replace_en_i;
    output [63:0] usr_rx5_data_o;
    output usr_rx5_pll_lock_o;
    input usr_rx5_pma_cdr_rst_i;
    input usr_rx5_pma_ckgen_rst_n_i;
    output usr_rx5_pma_loss_of_signal_o;
    input usr_rx5_pma_pll_rst_n_i;
    input usr_rx5_rst_n_i;
    input [3:0] usr_rx5_test_i;
    output [7:0] usr_rx5_test_o;
    output usr_tx0_busy_o;
    input [7:0] usr_tx0_ctrl_char_is_k_i;
    input [7:0] usr_tx0_ctrl_enc_en_i;
    input [7:0] usr_tx0_ctrl_end_of_frame_i;
    input [7:0] usr_tx0_ctrl_end_of_multiframe_i;
    input usr_tx0_ctrl_replace_en_i;
    input [7:0] usr_tx0_ctrl_scr_en_i;
    input [63:0] usr_tx0_data_i;
    input usr_tx0_pma_clk_en_i;
    input usr_tx0_rst_n_i;
    input [3:0] usr_tx0_test_i;
    output [3:0] usr_tx0_test_o;
    output usr_tx1_busy_o;
    input [7:0] usr_tx1_ctrl_char_is_k_i;
    input [7:0] usr_tx1_ctrl_enc_en_i;
    input [7:0] usr_tx1_ctrl_end_of_frame_i;
    input [7:0] usr_tx1_ctrl_end_of_multiframe_i;
    input usr_tx1_ctrl_replace_en_i;
    input [7:0] usr_tx1_ctrl_scr_en_i;
    input [63:0] usr_tx1_data_i;
    input usr_tx1_pma_clk_en_i;
    input usr_tx1_rst_n_i;
    input [3:0] usr_tx1_test_i;
    output [3:0] usr_tx1_test_o;
    output usr_tx2_busy_o;
    input [7:0] usr_tx2_ctrl_char_is_k_i;
    input [7:0] usr_tx2_ctrl_enc_en_i;
    input [7:0] usr_tx2_ctrl_end_of_frame_i;
    input [7:0] usr_tx2_ctrl_end_of_multiframe_i;
    input usr_tx2_ctrl_replace_en_i;
    input [7:0] usr_tx2_ctrl_scr_en_i;
    input [63:0] usr_tx2_data_i;
    input usr_tx2_pma_clk_en_i;
    input usr_tx2_rst_n_i;
    input [3:0] usr_tx2_test_i;
    output [3:0] usr_tx2_test_o;
    output usr_tx3_busy_o;
    input [7:0] usr_tx3_ctrl_char_is_k_i;
    input [7:0] usr_tx3_ctrl_enc_en_i;
    input [7:0] usr_tx3_ctrl_end_of_frame_i;
    input [7:0] usr_tx3_ctrl_end_of_multiframe_i;
    input usr_tx3_ctrl_replace_en_i;
    input [7:0] usr_tx3_ctrl_scr_en_i;
    input [63:0] usr_tx3_data_i;
    input usr_tx3_pma_clk_en_i;
    input usr_tx3_rst_n_i;
    input [3:0] usr_tx3_test_i;
    output [3:0] usr_tx3_test_o;
    output usr_tx4_busy_o;
    input [7:0] usr_tx4_ctrl_char_is_k_i;
    input [7:0] usr_tx4_ctrl_enc_en_i;
    input [7:0] usr_tx4_ctrl_end_of_frame_i;
    input [7:0] usr_tx4_ctrl_end_of_multiframe_i;
    input usr_tx4_ctrl_replace_en_i;
    input [7:0] usr_tx4_ctrl_scr_en_i;
    input [63:0] usr_tx4_data_i;
    input usr_tx4_pma_clk_en_i;
    input usr_tx4_rst_n_i;
    input [3:0] usr_tx4_test_i;
    output [3:0] usr_tx4_test_o;
    output usr_tx5_busy_o;
    input [7:0] usr_tx5_ctrl_char_is_k_i;
    input [7:0] usr_tx5_ctrl_enc_en_i;
    input [7:0] usr_tx5_ctrl_end_of_frame_i;
    input [7:0] usr_tx5_ctrl_end_of_multiframe_i;
    input usr_tx5_ctrl_replace_en_i;
    input [7:0] usr_tx5_ctrl_scr_en_i;
    input [63:0] usr_tx5_data_i;
    input usr_tx5_pma_clk_en_i;
    input usr_tx5_rst_n_i;
    input [3:0] usr_tx5_test_i;
    output [3:0] usr_tx5_test_o;
    parameter cfg_main_i = 34'b0000000000000000000000000000000000;
    parameter cfg_rx0_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx1_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx2_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx3_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx4_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_rx5_i = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter cfg_tx0_i = 0;
    parameter cfg_tx1_i = 0;
    parameter cfg_tx2_i = 0;
    parameter cfg_tx3_i = 0;
    parameter cfg_tx4_i = 0;
    parameter cfg_tx5_i = 0;
    parameter location = "";
endmodule

(* blackbox *)
module NX_HSSL_U_FULL(hssl_clk_user_tx_i, hssl_clk_user_rx_i, hssl_clk_ref_i, hssl_clock_o, hssl_rclock_o, usr_dyn_cfg_en_i, usr_dyn_cfg_calibration_cs_n_i, usr_dyn_cfg_we_n_i, usr_dyn_cfg_wdata_sel_i, usr_pll_pma_rst_n_i, usr_pll_pma_pwr_down_n_i, usr_main_rst_n_i, usr_pll_lock_o, usr_pll_pma_lock_analog_o, usr_pll_ckfb_lock_o, usr_calibrate_pma_out_o, usr_main_async_debug_ack_i, usr_main_async_debug_req_o, scan_en_i, usr_tx0_ctrl_replace_en_i, usr_tx0_rst_n_i
, usr_tx0_busy_o, usr_tx0_ctrl_invalid_k_o, usr_tx0_ctrl_driver_pwrdwn_n_i, usr_tx0_pma_clk_en_i, usr_tx0_pma_tx_clk_o, usr_rx0_ctrl_dscr_en_i, usr_rx0_ctrl_dec_en_i, usr_rx0_ctrl_align_en_i, usr_rx0_ctrl_align_sync_i, usr_rx0_ctrl_replace_en_i, usr_rx0_ctrl_el_buff_rst_i, usr_rx0_rst_n_i, usr_rx0_pma_rst_n_i, usr_rx0_pma_m_eye_rst_i, usr_rx0_pma_pwr_down_n_i, usr_rx0_ctrl_char_is_aligned_o, usr_rx0_ctrl_valid_realign_o, usr_rx0_busy_o, usr_rx0_pma_loss_of_signal_o, usr_rx0_pma_ll_fast_locked_o, usr_rx0_pma_ll_slow_locked_o
, usr_rx0_pma_pll_lock_o, usr_rx0_pma_pll_lock_track_o, usr_tx1_ctrl_replace_en_i, usr_tx1_rst_n_i, usr_tx1_busy_o, usr_tx1_ctrl_invalid_k_o, usr_tx1_ctrl_driver_pwrdwn_n_i, usr_tx1_pma_clk_en_i, usr_tx1_pma_tx_clk_o, usr_rx1_ctrl_dscr_en_i, usr_rx1_ctrl_dec_en_i, usr_rx1_ctrl_align_en_i, usr_rx1_ctrl_align_sync_i, usr_rx1_ctrl_replace_en_i, usr_rx1_ctrl_el_buff_rst_i, usr_rx1_rst_n_i, usr_rx1_pma_rst_n_i, usr_rx1_pma_m_eye_rst_i, usr_rx1_pma_pwr_down_n_i, usr_rx1_ctrl_char_is_aligned_o, usr_rx1_ctrl_valid_realign_o
, usr_rx1_busy_o, usr_rx1_pma_loss_of_signal_o, usr_rx1_pma_ll_fast_locked_o, usr_rx1_pma_ll_slow_locked_o, usr_rx1_pma_pll_lock_o, usr_rx1_pma_pll_lock_track_o, usr_tx2_ctrl_replace_en_i, usr_tx2_rst_n_i, usr_tx2_busy_o, usr_tx2_ctrl_invalid_k_o, usr_tx2_ctrl_driver_pwrdwn_n_i, usr_tx2_pma_clk_en_i, usr_tx2_pma_tx_clk_o, usr_rx2_ctrl_dscr_en_i, usr_rx2_ctrl_dec_en_i, usr_rx2_ctrl_align_en_i, usr_rx2_ctrl_align_sync_i, usr_rx2_ctrl_replace_en_i, usr_rx2_ctrl_el_buff_rst_i, usr_rx2_rst_n_i, usr_rx2_pma_rst_n_i
, usr_rx2_pma_m_eye_rst_i, usr_rx2_pma_pwr_down_n_i, usr_rx2_ctrl_char_is_aligned_o, usr_rx2_ctrl_valid_realign_o, usr_rx2_busy_o, usr_rx2_pma_loss_of_signal_o, usr_rx2_pma_ll_fast_locked_o, usr_rx2_pma_ll_slow_locked_o, usr_rx2_pma_pll_lock_o, usr_rx2_pma_pll_lock_track_o, usr_tx3_ctrl_replace_en_i, usr_tx3_rst_n_i, usr_tx3_busy_o, usr_tx3_ctrl_invalid_k_o, usr_tx3_ctrl_driver_pwrdwn_n_i, usr_tx3_pma_clk_en_i, usr_tx3_pma_tx_clk_o, usr_rx3_ctrl_dscr_en_i, usr_rx3_ctrl_dec_en_i, usr_rx3_ctrl_align_en_i, usr_rx3_ctrl_align_sync_i
, usr_rx3_ctrl_replace_en_i, usr_rx3_ctrl_el_buff_rst_i, usr_rx3_rst_n_i, usr_rx3_pma_rst_n_i, usr_rx3_pma_m_eye_rst_i, usr_rx3_pma_pwr_down_n_i, usr_rx3_ctrl_char_is_aligned_o, usr_rx3_ctrl_valid_realign_o, usr_rx3_busy_o, usr_rx3_pma_loss_of_signal_o, usr_rx3_pma_ll_fast_locked_o, usr_rx3_pma_ll_slow_locked_o, usr_rx3_pma_pll_lock_o, usr_rx3_pma_pll_lock_track_o, usr_tx0_ctrl_enc_en_i, usr_tx0_ctrl_char_is_k_i, usr_tx0_ctrl_scr_en_i, usr_tx0_ctrl_end_of_multiframe_i, usr_tx0_ctrl_end_of_frame_i, usr_tx0_data_i, usr_rx0_data_o
, usr_rx0_ctrl_ovs_bit_sel_i, usr_rx0_ctrl_char_is_comma_o, usr_rx0_ctrl_char_is_k_o, usr_rx0_ctrl_not_in_table_o, usr_rx0_ctrl_disp_err_o, usr_rx0_ctrl_char_is_a_o, usr_rx0_ctrl_char_is_f_o, usr_rx0_test_o, usr_tx1_ctrl_enc_en_i, usr_tx1_ctrl_char_is_k_i, usr_tx1_ctrl_scr_en_i, usr_tx1_ctrl_end_of_multiframe_i, usr_tx1_ctrl_end_of_frame_i, usr_tx1_data_i, usr_rx1_data_o, usr_rx1_ctrl_ovs_bit_sel_i, usr_rx1_ctrl_char_is_comma_o, usr_rx1_ctrl_char_is_k_o, usr_rx1_ctrl_not_in_table_o, usr_rx1_ctrl_disp_err_o, usr_rx1_ctrl_char_is_a_o
, usr_rx1_ctrl_char_is_f_o, usr_rx1_test_o, usr_tx2_ctrl_enc_en_i, usr_tx2_ctrl_char_is_k_i, usr_tx2_ctrl_scr_en_i, usr_tx2_ctrl_end_of_multiframe_i, usr_tx2_ctrl_end_of_frame_i, usr_tx2_data_i, usr_rx2_data_o, usr_rx2_ctrl_ovs_bit_sel_i, usr_rx2_ctrl_char_is_comma_o, usr_rx2_ctrl_char_is_k_o, usr_rx2_ctrl_not_in_table_o, usr_rx2_ctrl_disp_err_o, usr_rx2_ctrl_char_is_a_o, usr_rx2_ctrl_char_is_f_o, usr_rx2_test_o, usr_tx3_ctrl_enc_en_i, usr_tx3_ctrl_char_is_k_i, usr_tx3_ctrl_scr_en_i, usr_tx3_ctrl_end_of_multiframe_i
, usr_tx3_ctrl_end_of_frame_i, usr_tx3_data_i, usr_rx3_data_o, usr_rx3_ctrl_ovs_bit_sel_i, usr_rx3_ctrl_char_is_comma_o, usr_rx3_ctrl_char_is_k_o, usr_rx3_ctrl_not_in_table_o, usr_rx3_ctrl_disp_err_o, usr_rx3_ctrl_char_is_a_o, usr_rx3_ctrl_char_is_f_o, usr_rx3_test_o, usr_dyn_cfg_addr_i, usr_dyn_cfg_wdata_i, usr_main_async_debug_lane_sel_i, usr_main_rx_pma_ll_out_o, scan_in_i, scan_out_o, usr_rx0_ctrl_debug_sel_i, usr_rx1_ctrl_debug_sel_i, usr_rx2_ctrl_debug_sel_i, usr_rx3_ctrl_debug_sel_i
, usr_dyn_cfg_lane_cs_n_i);
    input hssl_clk_ref_i;
    input hssl_clk_user_rx_i;
    input hssl_clk_user_tx_i;
    output hssl_clock_o;
    output hssl_rclock_o;
    input scan_en_i;
    input [7:0] scan_in_i;
    output [7:0] scan_out_o;
    output usr_calibrate_pma_out_o;
    input [3:0] usr_dyn_cfg_addr_i;
    input usr_dyn_cfg_calibration_cs_n_i;
    input usr_dyn_cfg_en_i;
    input [3:0] usr_dyn_cfg_lane_cs_n_i;
    input [11:0] usr_dyn_cfg_wdata_i;
    input usr_dyn_cfg_wdata_sel_i;
    input usr_dyn_cfg_we_n_i;
    input usr_main_async_debug_ack_i;
    input [1:0] usr_main_async_debug_lane_sel_i;
    output usr_main_async_debug_req_o;
    input usr_main_rst_n_i;
    output [19:0] usr_main_rx_pma_ll_out_o;
    output usr_pll_ckfb_lock_o;
    output usr_pll_lock_o;
    output usr_pll_pma_lock_analog_o;
    input usr_pll_pma_pwr_down_n_i;
    input usr_pll_pma_rst_n_i;
    output usr_rx0_busy_o;
    input usr_rx0_ctrl_align_en_i;
    input usr_rx0_ctrl_align_sync_i;
    output [7:0] usr_rx0_ctrl_char_is_a_o;
    output usr_rx0_ctrl_char_is_aligned_o;
    output [7:0] usr_rx0_ctrl_char_is_comma_o;
    output [7:0] usr_rx0_ctrl_char_is_f_o;
    output [7:0] usr_rx0_ctrl_char_is_k_o;
    input [2:0] usr_rx0_ctrl_debug_sel_i;
    input usr_rx0_ctrl_dec_en_i;
    output [7:0] usr_rx0_ctrl_disp_err_o;
    input usr_rx0_ctrl_dscr_en_i;
    input usr_rx0_ctrl_el_buff_rst_i;
    output [7:0] usr_rx0_ctrl_not_in_table_o;
    input [1:0] usr_rx0_ctrl_ovs_bit_sel_i;
    input usr_rx0_ctrl_replace_en_i;
    output usr_rx0_ctrl_valid_realign_o;
    output [63:0] usr_rx0_data_o;
    output usr_rx0_pma_ll_fast_locked_o;
    output usr_rx0_pma_ll_slow_locked_o;
    output usr_rx0_pma_loss_of_signal_o;
    input usr_rx0_pma_m_eye_rst_i;
    output usr_rx0_pma_pll_lock_o;
    output usr_rx0_pma_pll_lock_track_o;
    input usr_rx0_pma_pwr_down_n_i;
    input usr_rx0_pma_rst_n_i;
    input usr_rx0_rst_n_i;
    output [7:0] usr_rx0_test_o;
    output usr_rx1_busy_o;
    input usr_rx1_ctrl_align_en_i;
    input usr_rx1_ctrl_align_sync_i;
    output [7:0] usr_rx1_ctrl_char_is_a_o;
    output usr_rx1_ctrl_char_is_aligned_o;
    output [7:0] usr_rx1_ctrl_char_is_comma_o;
    output [7:0] usr_rx1_ctrl_char_is_f_o;
    output [7:0] usr_rx1_ctrl_char_is_k_o;
    input [2:0] usr_rx1_ctrl_debug_sel_i;
    input usr_rx1_ctrl_dec_en_i;
    output [7:0] usr_rx1_ctrl_disp_err_o;
    input usr_rx1_ctrl_dscr_en_i;
    input usr_rx1_ctrl_el_buff_rst_i;
    output [7:0] usr_rx1_ctrl_not_in_table_o;
    input [1:0] usr_rx1_ctrl_ovs_bit_sel_i;
    input usr_rx1_ctrl_replace_en_i;
    output usr_rx1_ctrl_valid_realign_o;
    output [63:0] usr_rx1_data_o;
    output usr_rx1_pma_ll_fast_locked_o;
    output usr_rx1_pma_ll_slow_locked_o;
    output usr_rx1_pma_loss_of_signal_o;
    input usr_rx1_pma_m_eye_rst_i;
    output usr_rx1_pma_pll_lock_o;
    output usr_rx1_pma_pll_lock_track_o;
    input usr_rx1_pma_pwr_down_n_i;
    input usr_rx1_pma_rst_n_i;
    input usr_rx1_rst_n_i;
    output [7:0] usr_rx1_test_o;
    output usr_rx2_busy_o;
    input usr_rx2_ctrl_align_en_i;
    input usr_rx2_ctrl_align_sync_i;
    output [7:0] usr_rx2_ctrl_char_is_a_o;
    output usr_rx2_ctrl_char_is_aligned_o;
    output [7:0] usr_rx2_ctrl_char_is_comma_o;
    output [7:0] usr_rx2_ctrl_char_is_f_o;
    output [7:0] usr_rx2_ctrl_char_is_k_o;
    input [2:0] usr_rx2_ctrl_debug_sel_i;
    input usr_rx2_ctrl_dec_en_i;
    output [7:0] usr_rx2_ctrl_disp_err_o;
    input usr_rx2_ctrl_dscr_en_i;
    input usr_rx2_ctrl_el_buff_rst_i;
    output [7:0] usr_rx2_ctrl_not_in_table_o;
    input [1:0] usr_rx2_ctrl_ovs_bit_sel_i;
    input usr_rx2_ctrl_replace_en_i;
    output usr_rx2_ctrl_valid_realign_o;
    output [63:0] usr_rx2_data_o;
    output usr_rx2_pma_ll_fast_locked_o;
    output usr_rx2_pma_ll_slow_locked_o;
    output usr_rx2_pma_loss_of_signal_o;
    input usr_rx2_pma_m_eye_rst_i;
    output usr_rx2_pma_pll_lock_o;
    output usr_rx2_pma_pll_lock_track_o;
    input usr_rx2_pma_pwr_down_n_i;
    input usr_rx2_pma_rst_n_i;
    input usr_rx2_rst_n_i;
    output [7:0] usr_rx2_test_o;
    output usr_rx3_busy_o;
    input usr_rx3_ctrl_align_en_i;
    input usr_rx3_ctrl_align_sync_i;
    output [7:0] usr_rx3_ctrl_char_is_a_o;
    output usr_rx3_ctrl_char_is_aligned_o;
    output [7:0] usr_rx3_ctrl_char_is_comma_o;
    output [7:0] usr_rx3_ctrl_char_is_f_o;
    output [7:0] usr_rx3_ctrl_char_is_k_o;
    input [2:0] usr_rx3_ctrl_debug_sel_i;
    input usr_rx3_ctrl_dec_en_i;
    output [7:0] usr_rx3_ctrl_disp_err_o;
    input usr_rx3_ctrl_dscr_en_i;
    input usr_rx3_ctrl_el_buff_rst_i;
    output [7:0] usr_rx3_ctrl_not_in_table_o;
    input [1:0] usr_rx3_ctrl_ovs_bit_sel_i;
    input usr_rx3_ctrl_replace_en_i;
    output usr_rx3_ctrl_valid_realign_o;
    output [63:0] usr_rx3_data_o;
    output usr_rx3_pma_ll_fast_locked_o;
    output usr_rx3_pma_ll_slow_locked_o;
    output usr_rx3_pma_loss_of_signal_o;
    input usr_rx3_pma_m_eye_rst_i;
    output usr_rx3_pma_pll_lock_o;
    output usr_rx3_pma_pll_lock_track_o;
    input usr_rx3_pma_pwr_down_n_i;
    input usr_rx3_pma_rst_n_i;
    input usr_rx3_rst_n_i;
    output [7:0] usr_rx3_test_o;
    output usr_tx0_busy_o;
    input [7:0] usr_tx0_ctrl_char_is_k_i;
    input usr_tx0_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx0_ctrl_enc_en_i;
    input [7:0] usr_tx0_ctrl_end_of_frame_i;
    input [7:0] usr_tx0_ctrl_end_of_multiframe_i;
    output usr_tx0_ctrl_invalid_k_o;
    input usr_tx0_ctrl_replace_en_i;
    input [7:0] usr_tx0_ctrl_scr_en_i;
    input [63:0] usr_tx0_data_i;
    input usr_tx0_pma_clk_en_i;
    output usr_tx0_pma_tx_clk_o;
    input usr_tx0_rst_n_i;
    output usr_tx1_busy_o;
    input [7:0] usr_tx1_ctrl_char_is_k_i;
    input usr_tx1_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx1_ctrl_enc_en_i;
    input [7:0] usr_tx1_ctrl_end_of_frame_i;
    input [7:0] usr_tx1_ctrl_end_of_multiframe_i;
    output usr_tx1_ctrl_invalid_k_o;
    input usr_tx1_ctrl_replace_en_i;
    input [7:0] usr_tx1_ctrl_scr_en_i;
    input [63:0] usr_tx1_data_i;
    input usr_tx1_pma_clk_en_i;
    output usr_tx1_pma_tx_clk_o;
    input usr_tx1_rst_n_i;
    output usr_tx2_busy_o;
    input [7:0] usr_tx2_ctrl_char_is_k_i;
    input usr_tx2_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx2_ctrl_enc_en_i;
    input [7:0] usr_tx2_ctrl_end_of_frame_i;
    input [7:0] usr_tx2_ctrl_end_of_multiframe_i;
    output usr_tx2_ctrl_invalid_k_o;
    input usr_tx2_ctrl_replace_en_i;
    input [7:0] usr_tx2_ctrl_scr_en_i;
    input [63:0] usr_tx2_data_i;
    input usr_tx2_pma_clk_en_i;
    output usr_tx2_pma_tx_clk_o;
    input usr_tx2_rst_n_i;
    output usr_tx3_busy_o;
    input [7:0] usr_tx3_ctrl_char_is_k_i;
    input usr_tx3_ctrl_driver_pwrdwn_n_i;
    input [7:0] usr_tx3_ctrl_enc_en_i;
    input [7:0] usr_tx3_ctrl_end_of_frame_i;
    input [7:0] usr_tx3_ctrl_end_of_multiframe_i;
    output usr_tx3_ctrl_invalid_k_o;
    input usr_tx3_ctrl_replace_en_i;
    input [7:0] usr_tx3_ctrl_scr_en_i;
    input [63:0] usr_tx3_data_i;
    input usr_tx3_pma_clk_en_i;
    output usr_tx3_pma_tx_clk_o;
    input usr_tx3_rst_n_i;
    parameter cfg_dyn_all_rx_pma_m_eye_coarse_ena_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_dn_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_fine_ena_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_m_eye_step_i = 4'b0000;
    parameter cfg_dyn_all_rx_pma_m_eye_up_i = 1'b0;
    parameter cfg_dyn_all_rx_pma_threshold_1 = 5'b00000;
    parameter cfg_dyn_all_rx_pma_threshold_2 = 5'b00000;
    parameter cfg_dyn_all_rx_pma_trim_locked_i = 3'b000;
    parameter cfg_dyn_all_rx_pma_trim_mode_i = 2'b00;
    parameter cfg_dyn_all_rx_pma_trim_unlocked_i = 3'b000;
    parameter cfg_dyn_rx0_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx0_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx0_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx1_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx1_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx2_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx2_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_ctle_cap_p_i = 4'b0000;
    parameter cfg_dyn_rx3_pma_ctle_res_p_i = 4'b0000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap1_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap2_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap3_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_dfe_idac_tap4_n_i = 6'b000000;
    parameter cfg_dyn_rx3_pma_termination_cmd_i = 6'b000000;
    parameter cfg_dyn_tx0_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx0_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx0_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx0_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx0_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx0_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx0_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx0_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx0_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx0_pma_pre_sign_i = 1'b0;
    parameter cfg_dyn_tx1_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx1_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx1_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx1_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx1_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx1_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx1_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx1_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx1_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx1_pma_pre_sign_i = 1'b0;
    parameter cfg_dyn_tx2_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx2_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx2_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx2_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx2_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx2_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx2_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx2_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx2_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx2_pma_pre_sign_i = 1'b0;
    parameter cfg_dyn_tx3_pma_main_en_i = 6'b000000;
    parameter cfg_dyn_tx3_pma_main_sign_i = 1'b0;
    parameter cfg_dyn_tx3_pma_margin_input_i = 9'b000000000;
    parameter cfg_dyn_tx3_pma_margin_sel_i = 9'b000000000;
    parameter cfg_dyn_tx3_pma_post_en_i = 5'b00000;
    parameter cfg_dyn_tx3_pma_post_sel_i = 8'b00000000;
    parameter cfg_dyn_tx3_pma_post_sign_i = 1'b0;
    parameter cfg_dyn_tx3_pma_pre_en_i = 1'b0;
    parameter cfg_dyn_tx3_pma_pre_sel_i = 4'b0000;
    parameter cfg_dyn_tx3_pma_pre_sign_i = 1'b0;
    parameter cfg_main_clk_to_fabric_div_en_i = 1'b0;
    parameter cfg_main_clk_to_fabric_div_mode_i = 1'b0;
    parameter cfg_main_clk_to_fabric_sel_i = 1'b0;
    parameter cfg_main_rclk_to_fabric_sel_i = 2'b00;
    parameter cfg_main_use_only_usr_clock_i = 1'b0;
    parameter cfg_pcs_ovs_en_i = 1'b0;
    parameter cfg_pcs_ovs_mode_i = 1'b0;
    parameter cfg_pcs_pll_lock_ppm_i = 3'b000;
    parameter cfg_pcs_word_len_i = 2'b00;
    parameter cfg_pll_pma_ckref_ext_i = 1'b0;
    parameter cfg_pll_pma_cpump_i = 4'b0000;
    parameter cfg_pll_pma_divl_i = 2'b00;
    parameter cfg_pll_pma_divm_i = 1'b0;
    parameter cfg_pll_pma_divn_i = 2'b00;
    parameter cfg_pll_pma_gbx_en_i = 1'b0;
    parameter cfg_pll_pma_int_data_len_i = 1'b0;
    parameter cfg_pll_pma_lvds_en_i = 1'b0;
    parameter cfg_pll_pma_lvds_mux_i = 1'b0;
    parameter cfg_pll_pma_mux_ckref_i = 1'b0;
    parameter cfg_rx0_gearbox_en_i = 1'b0;
    parameter cfg_rx0_gearbox_mode_i = 1'b0;
    parameter cfg_rx0_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx0_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx0_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx0_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx0_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx0_pcs_debug_en_i = 1'b0;
    parameter cfg_rx0_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx0_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx0_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx0_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx0_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx0_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx0_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx0_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx0_pcs_loopback_i = 1'b0;
    parameter cfg_rx0_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx0_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx0_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx0_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx0_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx0_pcs_polarity_i = 1'b0;
    parameter cfg_rx0_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx0_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx0_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx0_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx0_pma_clk_pos_i = 1'b0;
    parameter cfg_rx0_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx0_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx0_pma_dco_divl_i = 2'b00;
    parameter cfg_rx0_pma_dco_divm_i = 1'b0;
    parameter cfg_rx0_pma_dco_divn_i = 2'b00;
    parameter cfg_rx0_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx0_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx0_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx0_pma_loopback_i = 1'b0;
    parameter cfg_rx0_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx0_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx0_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx0_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx0_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx0_pma_pll_divf_i = 2'b00;
    parameter cfg_rx0_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx0_pma_pll_divm_i = 2'b00;
    parameter cfg_rx0_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx0_pma_pll_divn_i = 1'b0;
    parameter cfg_rx1_gearbox_en_i = 1'b0;
    parameter cfg_rx1_gearbox_mode_i = 1'b0;
    parameter cfg_rx1_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx1_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx1_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx1_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx1_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx1_pcs_debug_en_i = 1'b0;
    parameter cfg_rx1_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx1_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx1_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx1_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx1_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx1_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx1_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx1_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx1_pcs_loopback_i = 1'b0;
    parameter cfg_rx1_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx1_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx1_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx1_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx1_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx1_pcs_polarity_i = 1'b0;
    parameter cfg_rx1_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx1_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx1_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx1_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx1_pma_clk_pos_i = 1'b0;
    parameter cfg_rx1_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx1_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx1_pma_dco_divl_i = 2'b00;
    parameter cfg_rx1_pma_dco_divm_i = 1'b0;
    parameter cfg_rx1_pma_dco_divn_i = 2'b00;
    parameter cfg_rx1_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx1_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx1_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx1_pma_loopback_i = 1'b0;
    parameter cfg_rx1_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx1_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx1_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx1_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx1_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx1_pma_pll_divf_i = 2'b00;
    parameter cfg_rx1_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx1_pma_pll_divm_i = 2'b00;
    parameter cfg_rx1_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx1_pma_pll_divn_i = 1'b0;
    parameter cfg_rx2_gearbox_en_i = 1'b0;
    parameter cfg_rx2_gearbox_mode_i = 1'b0;
    parameter cfg_rx2_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx2_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx2_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx2_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx2_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx2_pcs_debug_en_i = 1'b0;
    parameter cfg_rx2_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx2_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx2_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx2_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx2_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx2_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx2_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx2_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx2_pcs_loopback_i = 1'b0;
    parameter cfg_rx2_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx2_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx2_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx2_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx2_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx2_pcs_polarity_i = 1'b0;
    parameter cfg_rx2_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx2_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx2_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx2_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx2_pma_clk_pos_i = 1'b0;
    parameter cfg_rx2_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx2_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx2_pma_dco_divl_i = 2'b00;
    parameter cfg_rx2_pma_dco_divm_i = 1'b0;
    parameter cfg_rx2_pma_dco_divn_i = 2'b00;
    parameter cfg_rx2_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx2_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx2_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx2_pma_loopback_i = 1'b0;
    parameter cfg_rx2_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx2_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx2_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx2_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx2_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx2_pma_pll_divf_i = 2'b00;
    parameter cfg_rx2_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx2_pma_pll_divm_i = 2'b00;
    parameter cfg_rx2_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx2_pma_pll_divn_i = 1'b0;
    parameter cfg_rx3_gearbox_en_i = 1'b0;
    parameter cfg_rx3_gearbox_mode_i = 1'b0;
    parameter cfg_rx3_pcs_8b_dscr_sel_i = 1'b0;
    parameter cfg_rx3_pcs_align_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_buffers_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_buffers_use_cdc_i = 1'b0;
    parameter cfg_rx3_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_rx3_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_rx3_pcs_comma_mask_i = 10'b0000000000;
    parameter cfg_rx3_pcs_debug_en_i = 1'b0;
    parameter cfg_rx3_pcs_dec_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_dscr_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_el_buff_diff_bef_comp_i = 4'b0000;
    parameter cfg_rx3_pcs_el_buff_max_comp_i = 4'b0000;
    parameter cfg_rx3_pcs_el_buff_only_one_skp_i = 1'b0;
    parameter cfg_rx3_pcs_el_buff_skp_char_0_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_char_1_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_char_2_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_char_3_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_0_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_1_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_2_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_3_i = 9'b000000000;
    parameter cfg_rx3_pcs_el_buff_skp_header_size_i = 2'b00;
    parameter cfg_rx3_pcs_el_buff_skp_seq_size_i = 2'b00;
    parameter cfg_rx3_pcs_fsm_sel_i = 2'b00;
    parameter cfg_rx3_pcs_fsm_watchdog_en_i = 1'b0;
    parameter cfg_rx3_pcs_loopback_i = 1'b0;
    parameter cfg_rx3_pcs_m_comma_en_i = 1'b0;
    parameter cfg_rx3_pcs_m_comma_val_i = 10'b0000000000;
    parameter cfg_rx3_pcs_nb_comma_bef_realign_i = 2'b00;
    parameter cfg_rx3_pcs_p_comma_en_i = 1'b0;
    parameter cfg_rx3_pcs_p_comma_val_i = 10'b0000000000;
    parameter cfg_rx3_pcs_polarity_i = 1'b0;
    parameter cfg_rx3_pcs_protocol_size_i = 1'b0;
    parameter cfg_rx3_pcs_replace_bypass_i = 1'b0;
    parameter cfg_rx3_pcs_sync_supported_i = 1'b0;
    parameter cfg_rx3_pma_cdr_cp_i = 4'b0000;
    parameter cfg_rx3_pma_clk_pos_i = 1'b0;
    parameter cfg_rx3_pma_coarse_ppm_i = 3'b000;
    parameter cfg_rx3_pma_ctrl_term_i = 6'b000000;
    parameter cfg_rx3_pma_dco_divl_i = 2'b00;
    parameter cfg_rx3_pma_dco_divm_i = 1'b0;
    parameter cfg_rx3_pma_dco_divn_i = 2'b00;
    parameter cfg_rx3_pma_dco_reg_res_i = 2'b00;
    parameter cfg_rx3_pma_dco_vref_sel_i = 1'b0;
    parameter cfg_rx3_pma_fine_ppm_i = 3'b000;
    parameter cfg_rx3_pma_loopback_i = 1'b0;
    parameter cfg_rx3_pma_m_eye_ppm_i = 3'b000;
    parameter cfg_rx3_pma_peak_detect_cmd_i = 2'b00;
    parameter cfg_rx3_pma_peak_detect_on_i = 1'b0;
    parameter cfg_rx3_pma_pll_cpump_n_i = 3'b000;
    parameter cfg_rx3_pma_pll_divf_en_n_i = 1'b0;
    parameter cfg_rx3_pma_pll_divf_i = 2'b00;
    parameter cfg_rx3_pma_pll_divm_en_n_i = 1'b0;
    parameter cfg_rx3_pma_pll_divm_i = 2'b00;
    parameter cfg_rx3_pma_pll_divn_en_n_i = 1'b0;
    parameter cfg_rx3_pma_pll_divn_i = 1'b0;
    parameter cfg_test_mode_i = 2'b00;
    parameter cfg_tx0_gearbox_en_i = 1'b0;
    parameter cfg_tx0_gearbox_mode_i = 1'b0;
    parameter cfg_tx0_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx0_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx0_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx0_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx0_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx0_pcs_loopback_i = 1'b0;
    parameter cfg_tx0_pcs_polarity_i = 1'b0;
    parameter cfg_tx0_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx0_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx0_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx0_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx0_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx0_pma_clk_pos_i = 1'b0;
    parameter cfg_tx0_pma_loopback_i = 1'b0;
    parameter cfg_tx1_gearbox_en_i = 1'b0;
    parameter cfg_tx1_gearbox_mode_i = 1'b0;
    parameter cfg_tx1_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx1_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx1_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx1_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx1_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx1_pcs_loopback_i = 1'b0;
    parameter cfg_tx1_pcs_polarity_i = 1'b0;
    parameter cfg_tx1_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx1_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx1_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx1_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx1_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx1_pma_clk_pos_i = 1'b0;
    parameter cfg_tx1_pma_loopback_i = 1'b0;
    parameter cfg_tx2_gearbox_en_i = 1'b0;
    parameter cfg_tx2_gearbox_mode_i = 1'b0;
    parameter cfg_tx2_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx2_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx2_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx2_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx2_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx2_pcs_loopback_i = 1'b0;
    parameter cfg_tx2_pcs_polarity_i = 1'b0;
    parameter cfg_tx2_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx2_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx2_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx2_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx2_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx2_pma_clk_pos_i = 1'b0;
    parameter cfg_tx2_pma_loopback_i = 1'b0;
    parameter cfg_tx3_gearbox_en_i = 1'b0;
    parameter cfg_tx3_gearbox_mode_i = 1'b0;
    parameter cfg_tx3_pcs_8b_scr_sel_i = 1'b0;
    parameter cfg_tx3_pcs_bypass_pma_cdc_i = 1'b0;
    parameter cfg_tx3_pcs_bypass_usr_cdc_i = 1'b0;
    parameter cfg_tx3_pcs_enc_bypass_i = 1'b0;
    parameter cfg_tx3_pcs_esistream_fsm_en_i = 1'b0;
    parameter cfg_tx3_pcs_loopback_i = 1'b0;
    parameter cfg_tx3_pcs_polarity_i = 1'b0;
    parameter cfg_tx3_pcs_protocol_size_i = 1'b0;
    parameter cfg_tx3_pcs_replace_bypass_i = 1'b0;
    parameter cfg_tx3_pcs_scr_bypass_i = 1'b0;
    parameter cfg_tx3_pcs_scr_init_i = 17'b00000000000000000;
    parameter cfg_tx3_pcs_sync_supported_i = 1'b0;
    parameter cfg_tx3_pma_clk_pos_i = 1'b0;
    parameter cfg_tx3_pma_loopback_i = 1'b0;
    parameter location = "";
    parameter rx_usrclk_use_pcs_clk_2 = 1'b0;
    parameter tx_usrclk_use_pcs_clk_2 = 1'b0;
endmodule

(* blackbox *)
module NX_IOB(I, C, T, O, IO);
    input C;
    input I;
    inout IO;
    output O;
    input T;
    parameter differential = "";
    parameter drive = "";
    parameter dynDrive = "";
    parameter dynInput = "";
    parameter dynTerm = "";
    parameter extra = 3;
    parameter inputDelayLine = "";
    parameter inputDelayOn = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter outputDelayOn = "";
    parameter slewRate = "";
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_IOB_I(C, T, IO, O);
    input C;
    input IO;
    output O;
    input T;
    parameter differential = "";
    parameter drive = "";
    parameter dynDrive = "";
    parameter dynInput = "";
    parameter dynTerm = "";
    parameter extra = 1;
    parameter inputDelayLine = "";
    parameter inputDelayOn = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter outputDelayOn = "";
    parameter slewRate = "";
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_IOB_O(I, C, T, IO);
    input C;
    input I;
    output IO;
    input T;
    parameter differential = "";
    parameter drive = "";
    parameter dynDrive = "";
    parameter dynInput = "";
    parameter dynTerm = "";
    parameter extra = 2;
    parameter inputDelayLine = "";
    parameter inputDelayOn = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter outputDelayOn = "";
    parameter slewRate = "";
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_IOM(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, CCK, DCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1
, C2RW2, C2RW3, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FZ, DC, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3, DRA4
, DRA5, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1, CAP2, CAP3
, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, SPI1, SPI2, SPI3, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1, DRO2, DRO3
, DRO4, DRO5, DRO6, CAL, P1CI1, P1CL, P1CR, P1CO, P1CTI, P1CTO, P1EI1, P1EI2, P1EI3, P1EI4, P1EI5, P1EL, P1ER, P1EO, P1RI, P1RL, P1RR
, P1RO1, P1RO2, P1RO3, P1RO4, P1RO5, P2CI1, P2CL, P2CR, P2CO, P2CTI, P2CTO, P2EI1, P2EI2, P2EI3, P2EI4, P2EI5, P2EL, P2ER, P2EO, P2RI, P2RL
, P2RR, P2RO1, P2RO2, P2RO3, P2RO4, P2RO5, P3CI1, P3CL, P3CR, P3CO, P3CTI, P3CTO, P3EI1, P3EI2, P3EI3, P3EI4, P3EI5, P3EL, P3ER, P3EO, P3RI
, P3RL, P3RR, P3RO1, P3RO2, P3RO3, P3RO4, P3RO5, P4CI1, P4CL, P4CR, P4CO, P4CTI, P4CTO, P4EI1, P4EI2, P4EI3, P4EI4, P4EI5, P4EL, P4ER, P4EO
, P4RI, P4RL, P4RR, P4RO1, P4RO2, P4RO3, P4RO4, P4RO5, P5CI1, P5CI2, P5CI3, P5CI4, P5CI5, P5CL, P5CR, P5CO, P5CTI, P5CTO, P5EI1, P5EI2, P5EI3
, P5EI4, P5EI5, P5EL, P5ER, P5EO, P5RI, P5RL, P5RR, P5RO1, P5RO2, P5RO3, P5RO4, P5RO5, P6CI1, P6CL, P6CR, P6CO, P6CTI, P6CTO, P6EI1, P6EI2
, P6EI3, P6EI4, P6EI5, P6EL, P6ER, P6EO, P6RI, P6RL, P6RR, P6RO1, P6RO2, P6RO3, P6RO4, P6RO5, P7CI1, P7CL, P7CR, P7CO, P7CTI, P7CTO, P7EI1
, P7EI2, P7EI3, P7EI4, P7EI5, P7EL, P7ER, P7EO, P7RI, P7RL, P7RR, P7RO1, P7RO2, P7RO3, P7RO4, P7RO5, P8CI1, P8CL, P8CR, P8CO, P8CTI, P8CTO
, P8EI1, P8EI2, P8EI3, P8EI4, P8EI5, P8EL, P8ER, P8EO, P8RI, P8RL, P8RR, P8RO1, P8RO2, P8RO3, P8RO4, P8RO5, P9CI1, P9CL, P9CR, P9CO, P9CTI
, P9CTO, P9EI1, P9EI2, P9EI3, P9EI4, P9EI5, P9EL, P9ER, P9EO, P9RI, P9RL, P9RR, P9RO1, P9RO2, P9RO3, P9RO4, P9RO5, P10CI1, P10CL, P10CR, P10CO
, P10CTI, P10CTO, P10EI1, P10EI2, P10EI3, P10EI4, P10EI5, P10EL, P10ER, P10EO, P10RI, P10RL, P10RR, P10RO1, P10RO2, P10RO3, P10RO4, P10RO5, P11CI1, P11CL, P11CR
, P11CO, P11CTI, P11CTO, P11EI1, P11EI2, P11EI3, P11EI4, P11EI5, P11EL, P11ER, P11EO, P11RI, P11RL, P11RR, P11RO1, P11RO2, P11RO3, P11RO4, P11RO5, P12CI1, P12CL
, P12CR, P12CO, P12CTI, P12CTO, P12EI1, P12EI2, P12EI3, P12EI4, P12EI5, P12EL, P12ER, P12EO, P12RI, P12RL, P12RR, P12RO1, P12RO2, P12RO3, P12RO4, P12RO5, P13CI1
, P13CL, P13CR, P13CO, P13CTI, P13CTO, P13EI1, P13EI2, P13EI3, P13EI4, P13EI5, P13EL, P13ER, P13EO, P13RI, P13RL, P13RR, P13RO1, P13RO2, P13RO3, P13RO4, P13RO5
, P14CI1, P14CL, P14CR, P14CO, P14CTI, P14CTO, P14EI1, P14EI2, P14EI3, P14EI4, P14EI5, P14EL, P14ER, P14EO, P14RI, P14RL, P14RR, P14RO1, P14RO2, P14RO3, P14RO4
, P14RO5, P15CI1, P15CL, P15CR, P15CO, P15CTI, P15CTO, P15EI1, P15EI2, P15EI3, P15EI4, P15EI5, P15EL, P15ER, P15EO, P15RI, P15RL, P15RR, P15RO1, P15RO2, P15RO3
, P15RO4, P15RO5, P16CI1, P16CL, P16CR, P16CO, P16CTI, P16CTO, P16EI1, P16EI2, P16EI3, P16EI4, P16EI5, P16EL, P16ER, P16EO, P16RI, P16RL, P16RR, P16RO1, P16RO2
, P16RO3, P16RO4, P16RO5, P17CI1, P17CL, P17CR, P17CO, P17CTI, P17CTO, P17EI1, P17EI2, P17EI3, P17EI4, P17EI5, P17EL, P17ER, P17EO, P17RI, P17RL, P17RR, P17RO1
, P17RO2, P17RO3, P17RO4, P17RO5, P18CI1, P18CL, P18CR, P18CO, P18CTI, P18CTO, P18EI1, P18EI2, P18EI3, P18EI4, P18EI5, P18EL, P18ER, P18EO, P18RI, P18RL, P18RR
, P18RO1, P18RO2, P18RO3, P18RO4, P18RO5, P19CI1, P19CL, P19CR, P19CO, P19CTI, P19CTO, P19EI1, P19EI2, P19EI3, P19EI4, P19EI5, P19EL, P19ER, P19EO, P19RI, P19RL
, P19RR, P19RO1, P19RO2, P19RO3, P19RO4, P19RO5, P20CI1, P20CL, P20CR, P20CO, P20CTI, P20CTO, P20EI1, P20EI2, P20EI3, P20EI4, P20EI5, P20EL, P20ER, P20EO, P20RI
, P20RL, P20RR, P20RO1, P20RO2, P20RO3, P20RO4, P20RO5, P21CI1, P21CL, P21CR, P21CO, P21CTI, P21CTO, P21EI1, P21EI2, P21EI3, P21EI4, P21EI5, P21EL, P21ER, P21EO
, P21RI, P21RL, P21RR, P21RO1, P21RO2, P21RO3, P21RO4, P21RO5, P22CI1, P22CL, P22CR, P22CO, P22CTI, P22CTO, P22EI1, P22EI2, P22EI3, P22EI4, P22EI5, P22EL, P22ER
, P22EO, P22RI, P22RL, P22RR, P22RO1, P22RO2, P22RO3, P22RO4, P22RO5, P23CI1, P23CL, P23CR, P23CO, P23CTI, P23CTO, P23EI1, P23EI2, P23EI3, P23EI4, P23EI5, P23EL
, P23ER, P23EO, P23RI, P23RL, P23RR, P23RO1, P23RO2, P23RO3, P23RO4, P23RO5, P24CI1, P24CL, P24CR, P24CO, P24CTI, P24CTO, P24EI1, P24EI2, P24EI3, P24EI4, P24EI5
, P24EL, P24ER, P24EO, P24RI, P24RL, P24RR, P24RO1, P24RO2, P24RO3, P24RO4, P24RO5, P25CI1, P25CI2, P25CI3, P25CI4, P25CI5, P25CL, P25CR, P25CO, P25CTI, P25CTO
, P25EI1, P25EI2, P25EI3, P25EI4, P25EI5, P25EL, P25ER, P25EO, P25RI, P25RL, P25RR, P25RO1, P25RO2, P25RO3, P25RO4, P25RO5, P26CI1, P26CL, P26CR, P26CO, P26CTI
, P26CTO, P26EI1, P26EI2, P26EI3, P26EI4, P26EI5, P26EL, P26ER, P26EO, P26RI, P26RL, P26RR, P26RO1, P26RO2, P26RO3, P26RO4, P26RO5, P27CI1, P27CL, P27CR, P27CO
, P27CTI, P27CTO, P27EI1, P27EI2, P27EI3, P27EI4, P27EI5, P27EL, P27ER, P27EO, P27RI, P27RL, P27RR, P27RO1, P27RO2, P27RO3, P27RO4, P27RO5, P28CI1, P28CL, P28CR
, P28CO, P28CTI, P28CTO, P28EI1, P28EI2, P28EI3, P28EI4, P28EI5, P28EL, P28ER, P28EO, P28RI, P28RL, P28RR, P28RO1, P28RO2, P28RO3, P28RO4, P28RO5, P29CI1, P29CL
, P29CR, P29CO, P29CTI, P29CTO, P29EI1, P29EI2, P29EI3, P29EI4, P29EI5, P29EL, P29ER, P29EO, P29RI, P29RL, P29RR, P29RO1, P29RO2, P29RO3, P29RO4, P29RO5, P30CI1
, P30CL, P30CR, P30CO, P30CTI, P30CTO, P30EI1, P30EI2, P30EI3, P30EI4, P30EI5, P30EL, P30ER, P30EO, P30RI, P30RL, P30RR, P30RO1, P30RO2, P30RO3, P30RO4, P30RO5
);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    output FLD;
    output FLG;
    input FZ;
    input P10CI1;
    input P10CL;
    output P10CO;
    input P10CR;
    input P10CTI;
    output P10CTO;
    input P10EI1;
    input P10EI2;
    input P10EI3;
    input P10EI4;
    input P10EI5;
    input P10EL;
    output P10EO;
    input P10ER;
    input P10RI;
    input P10RL;
    output P10RO1;
    output P10RO2;
    output P10RO3;
    output P10RO4;
    output P10RO5;
    input P10RR;
    input P11CI1;
    input P11CL;
    output P11CO;
    input P11CR;
    input P11CTI;
    output P11CTO;
    input P11EI1;
    input P11EI2;
    input P11EI3;
    input P11EI4;
    input P11EI5;
    input P11EL;
    output P11EO;
    input P11ER;
    input P11RI;
    input P11RL;
    output P11RO1;
    output P11RO2;
    output P11RO3;
    output P11RO4;
    output P11RO5;
    input P11RR;
    input P12CI1;
    input P12CL;
    output P12CO;
    input P12CR;
    input P12CTI;
    output P12CTO;
    input P12EI1;
    input P12EI2;
    input P12EI3;
    input P12EI4;
    input P12EI5;
    input P12EL;
    output P12EO;
    input P12ER;
    input P12RI;
    input P12RL;
    output P12RO1;
    output P12RO2;
    output P12RO3;
    output P12RO4;
    output P12RO5;
    input P12RR;
    input P13CI1;
    input P13CL;
    output P13CO;
    input P13CR;
    input P13CTI;
    output P13CTO;
    input P13EI1;
    input P13EI2;
    input P13EI3;
    input P13EI4;
    input P13EI5;
    input P13EL;
    output P13EO;
    input P13ER;
    input P13RI;
    input P13RL;
    output P13RO1;
    output P13RO2;
    output P13RO3;
    output P13RO4;
    output P13RO5;
    input P13RR;
    input P14CI1;
    input P14CL;
    output P14CO;
    input P14CR;
    input P14CTI;
    output P14CTO;
    input P14EI1;
    input P14EI2;
    input P14EI3;
    input P14EI4;
    input P14EI5;
    input P14EL;
    output P14EO;
    input P14ER;
    input P14RI;
    input P14RL;
    output P14RO1;
    output P14RO2;
    output P14RO3;
    output P14RO4;
    output P14RO5;
    input P14RR;
    input P15CI1;
    input P15CL;
    output P15CO;
    input P15CR;
    input P15CTI;
    output P15CTO;
    input P15EI1;
    input P15EI2;
    input P15EI3;
    input P15EI4;
    input P15EI5;
    input P15EL;
    output P15EO;
    input P15ER;
    input P15RI;
    input P15RL;
    output P15RO1;
    output P15RO2;
    output P15RO3;
    output P15RO4;
    output P15RO5;
    input P15RR;
    input P16CI1;
    input P16CL;
    output P16CO;
    input P16CR;
    input P16CTI;
    output P16CTO;
    input P16EI1;
    input P16EI2;
    input P16EI3;
    input P16EI4;
    input P16EI5;
    input P16EL;
    output P16EO;
    input P16ER;
    input P16RI;
    input P16RL;
    output P16RO1;
    output P16RO2;
    output P16RO3;
    output P16RO4;
    output P16RO5;
    input P16RR;
    input P17CI1;
    input P17CL;
    output P17CO;
    input P17CR;
    input P17CTI;
    output P17CTO;
    input P17EI1;
    input P17EI2;
    input P17EI3;
    input P17EI4;
    input P17EI5;
    input P17EL;
    output P17EO;
    input P17ER;
    input P17RI;
    input P17RL;
    output P17RO1;
    output P17RO2;
    output P17RO3;
    output P17RO4;
    output P17RO5;
    input P17RR;
    input P18CI1;
    input P18CL;
    output P18CO;
    input P18CR;
    input P18CTI;
    output P18CTO;
    input P18EI1;
    input P18EI2;
    input P18EI3;
    input P18EI4;
    input P18EI5;
    input P18EL;
    output P18EO;
    input P18ER;
    input P18RI;
    input P18RL;
    output P18RO1;
    output P18RO2;
    output P18RO3;
    output P18RO4;
    output P18RO5;
    input P18RR;
    input P19CI1;
    input P19CL;
    output P19CO;
    input P19CR;
    input P19CTI;
    output P19CTO;
    input P19EI1;
    input P19EI2;
    input P19EI3;
    input P19EI4;
    input P19EI5;
    input P19EL;
    output P19EO;
    input P19ER;
    input P19RI;
    input P19RL;
    output P19RO1;
    output P19RO2;
    output P19RO3;
    output P19RO4;
    output P19RO5;
    input P19RR;
    input P1CI1;
    input P1CL;
    output P1CO;
    input P1CR;
    input P1CTI;
    output P1CTO;
    input P1EI1;
    input P1EI2;
    input P1EI3;
    input P1EI4;
    input P1EI5;
    input P1EL;
    output P1EO;
    input P1ER;
    input P1RI;
    input P1RL;
    output P1RO1;
    output P1RO2;
    output P1RO3;
    output P1RO4;
    output P1RO5;
    input P1RR;
    input P20CI1;
    input P20CL;
    output P20CO;
    input P20CR;
    input P20CTI;
    output P20CTO;
    input P20EI1;
    input P20EI2;
    input P20EI3;
    input P20EI4;
    input P20EI5;
    input P20EL;
    output P20EO;
    input P20ER;
    input P20RI;
    input P20RL;
    output P20RO1;
    output P20RO2;
    output P20RO3;
    output P20RO4;
    output P20RO5;
    input P20RR;
    input P21CI1;
    input P21CL;
    output P21CO;
    input P21CR;
    input P21CTI;
    output P21CTO;
    input P21EI1;
    input P21EI2;
    input P21EI3;
    input P21EI4;
    input P21EI5;
    input P21EL;
    output P21EO;
    input P21ER;
    input P21RI;
    input P21RL;
    output P21RO1;
    output P21RO2;
    output P21RO3;
    output P21RO4;
    output P21RO5;
    input P21RR;
    input P22CI1;
    input P22CL;
    output P22CO;
    input P22CR;
    input P22CTI;
    output P22CTO;
    input P22EI1;
    input P22EI2;
    input P22EI3;
    input P22EI4;
    input P22EI5;
    input P22EL;
    output P22EO;
    input P22ER;
    input P22RI;
    input P22RL;
    output P22RO1;
    output P22RO2;
    output P22RO3;
    output P22RO4;
    output P22RO5;
    input P22RR;
    input P23CI1;
    input P23CL;
    output P23CO;
    input P23CR;
    input P23CTI;
    output P23CTO;
    input P23EI1;
    input P23EI2;
    input P23EI3;
    input P23EI4;
    input P23EI5;
    input P23EL;
    output P23EO;
    input P23ER;
    input P23RI;
    input P23RL;
    output P23RO1;
    output P23RO2;
    output P23RO3;
    output P23RO4;
    output P23RO5;
    input P23RR;
    input P24CI1;
    input P24CL;
    output P24CO;
    input P24CR;
    input P24CTI;
    output P24CTO;
    input P24EI1;
    input P24EI2;
    input P24EI3;
    input P24EI4;
    input P24EI5;
    input P24EL;
    output P24EO;
    input P24ER;
    input P24RI;
    input P24RL;
    output P24RO1;
    output P24RO2;
    output P24RO3;
    output P24RO4;
    output P24RO5;
    input P24RR;
    input P25CI1;
    input P25CI2;
    input P25CI3;
    input P25CI4;
    input P25CI5;
    input P25CL;
    output P25CO;
    input P25CR;
    input P25CTI;
    output P25CTO;
    input P25EI1;
    input P25EI2;
    input P25EI3;
    input P25EI4;
    input P25EI5;
    input P25EL;
    output P25EO;
    input P25ER;
    input P25RI;
    input P25RL;
    output P25RO1;
    output P25RO2;
    output P25RO3;
    output P25RO4;
    output P25RO5;
    input P25RR;
    input P26CI1;
    input P26CL;
    output P26CO;
    input P26CR;
    input P26CTI;
    output P26CTO;
    input P26EI1;
    input P26EI2;
    input P26EI3;
    input P26EI4;
    input P26EI5;
    input P26EL;
    output P26EO;
    input P26ER;
    input P26RI;
    input P26RL;
    output P26RO1;
    output P26RO2;
    output P26RO3;
    output P26RO4;
    output P26RO5;
    input P26RR;
    input P27CI1;
    input P27CL;
    output P27CO;
    input P27CR;
    input P27CTI;
    output P27CTO;
    input P27EI1;
    input P27EI2;
    input P27EI3;
    input P27EI4;
    input P27EI5;
    input P27EL;
    output P27EO;
    input P27ER;
    input P27RI;
    input P27RL;
    output P27RO1;
    output P27RO2;
    output P27RO3;
    output P27RO4;
    output P27RO5;
    input P27RR;
    input P28CI1;
    input P28CL;
    output P28CO;
    input P28CR;
    input P28CTI;
    output P28CTO;
    input P28EI1;
    input P28EI2;
    input P28EI3;
    input P28EI4;
    input P28EI5;
    input P28EL;
    output P28EO;
    input P28ER;
    input P28RI;
    input P28RL;
    output P28RO1;
    output P28RO2;
    output P28RO3;
    output P28RO4;
    output P28RO5;
    input P28RR;
    input P29CI1;
    input P29CL;
    output P29CO;
    input P29CR;
    input P29CTI;
    output P29CTO;
    input P29EI1;
    input P29EI2;
    input P29EI3;
    input P29EI4;
    input P29EI5;
    input P29EL;
    output P29EO;
    input P29ER;
    input P29RI;
    input P29RL;
    output P29RO1;
    output P29RO2;
    output P29RO3;
    output P29RO4;
    output P29RO5;
    input P29RR;
    input P2CI1;
    input P2CL;
    output P2CO;
    input P2CR;
    input P2CTI;
    output P2CTO;
    input P2EI1;
    input P2EI2;
    input P2EI3;
    input P2EI4;
    input P2EI5;
    input P2EL;
    output P2EO;
    input P2ER;
    input P2RI;
    input P2RL;
    output P2RO1;
    output P2RO2;
    output P2RO3;
    output P2RO4;
    output P2RO5;
    input P2RR;
    input P30CI1;
    input P30CL;
    output P30CO;
    input P30CR;
    input P30CTI;
    output P30CTO;
    input P30EI1;
    input P30EI2;
    input P30EI3;
    input P30EI4;
    input P30EI5;
    input P30EL;
    output P30EO;
    input P30ER;
    input P30RI;
    input P30RL;
    output P30RO1;
    output P30RO2;
    output P30RO3;
    output P30RO4;
    output P30RO5;
    input P30RR;
    input P3CI1;
    input P3CL;
    output P3CO;
    input P3CR;
    input P3CTI;
    output P3CTO;
    input P3EI1;
    input P3EI2;
    input P3EI3;
    input P3EI4;
    input P3EI5;
    input P3EL;
    output P3EO;
    input P3ER;
    input P3RI;
    input P3RL;
    output P3RO1;
    output P3RO2;
    output P3RO3;
    output P3RO4;
    output P3RO5;
    input P3RR;
    input P4CI1;
    input P4CL;
    output P4CO;
    input P4CR;
    input P4CTI;
    output P4CTO;
    input P4EI1;
    input P4EI2;
    input P4EI3;
    input P4EI4;
    input P4EI5;
    input P4EL;
    output P4EO;
    input P4ER;
    input P4RI;
    input P4RL;
    output P4RO1;
    output P4RO2;
    output P4RO3;
    output P4RO4;
    output P4RO5;
    input P4RR;
    input P5CI1;
    input P5CI2;
    input P5CI3;
    input P5CI4;
    input P5CI5;
    input P5CL;
    output P5CO;
    input P5CR;
    input P5CTI;
    output P5CTO;
    input P5EI1;
    input P5EI2;
    input P5EI3;
    input P5EI4;
    input P5EI5;
    input P5EL;
    output P5EO;
    input P5ER;
    input P5RI;
    input P5RL;
    output P5RO1;
    output P5RO2;
    output P5RO3;
    output P5RO4;
    output P5RO5;
    input P5RR;
    input P6CI1;
    input P6CL;
    output P6CO;
    input P6CR;
    input P6CTI;
    output P6CTO;
    input P6EI1;
    input P6EI2;
    input P6EI3;
    input P6EI4;
    input P6EI5;
    input P6EL;
    output P6EO;
    input P6ER;
    input P6RI;
    input P6RL;
    output P6RO1;
    output P6RO2;
    output P6RO3;
    output P6RO4;
    output P6RO5;
    input P6RR;
    input P7CI1;
    input P7CL;
    output P7CO;
    input P7CR;
    input P7CTI;
    output P7CTO;
    input P7EI1;
    input P7EI2;
    input P7EI3;
    input P7EI4;
    input P7EI5;
    input P7EL;
    output P7EO;
    input P7ER;
    input P7RI;
    input P7RL;
    output P7RO1;
    output P7RO2;
    output P7RO3;
    output P7RO4;
    output P7RO5;
    input P7RR;
    input P8CI1;
    input P8CL;
    output P8CO;
    input P8CR;
    input P8CTI;
    output P8CTO;
    input P8EI1;
    input P8EI2;
    input P8EI3;
    input P8EI4;
    input P8EI5;
    input P8EL;
    output P8EO;
    input P8ER;
    input P8RI;
    input P8RL;
    output P8RO1;
    output P8RO2;
    output P8RO3;
    output P8RO4;
    output P8RO5;
    input P8RR;
    input P9CI1;
    input P9CL;
    output P9CO;
    input P9CR;
    input P9CTI;
    output P9CTO;
    input P9EI1;
    input P9EI2;
    input P9EI3;
    input P9EI4;
    input P9EI5;
    input P9EL;
    output P9EO;
    input P9ER;
    input P9RI;
    input P9RL;
    output P9RO1;
    output P9RO2;
    output P9RO3;
    output P9RO4;
    output P9RO5;
    input P9RR;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input SPI1;
    input SPI2;
    input SPI3;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter mode_io_cal = 1'b0;
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter pads_dict = "";
    parameter pads_path = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_BIN2GRP(GS, DS, GVON, GVIN, GVDN, PA, LA);
    input [1:0] DS;
    input GS;
    output [2:0] GVDN;
    output [2:0] GVIN;
    output [2:0] GVON;
    input [5:0] LA;
    output [3:0] PA;
endmodule

(* blackbox *)
module NX_IOM_CONTROL(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1, C2RW2, C2RW3
, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, CCK, DCK, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, SPI1, SPI2, SPI3, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1
, DRO2, DRO3, DRO4, DRO5, DRO6, CAL, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16
, LINK17, LINK18, LINK19, LINK20, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input SPI1;
    input SPI2;
    input SPI3;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter inv_di_fclk1 = 1'b0;
    parameter inv_di_fclk2 = 1'b0;
    parameter latency1 = 1'b0;
    parameter latency2 = 1'b0;
    parameter location = "";
    parameter mode_cpath = "";
    parameter mode_epath = "";
    parameter mode_io_cal = 1'b0;
    parameter mode_rpath = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_tpath = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_CONTROL_L(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1, C2RW2, C2RW3
, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, CCK, DCK, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1, DRO2, DRO3, DRO4
, DRO5, DRO6, CAL, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16, LINK17, LINK18, LINK19
, LINK20, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter inv_di_fclk1 = 1'b0;
    parameter inv_di_fclk2 = 1'b0;
    parameter latency1 = 1'b0;
    parameter latency2 = 1'b0;
    parameter location = "";
    parameter mode_cpath = "";
    parameter mode_epath = "";
    parameter mode_io_cal = 1'b0;
    parameter mode_rpath = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_tpath = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_CONTROL_M(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1, C2RW2, C2RW3
, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, CCK, DCK, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, SPI1, SPI2, SPI3, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1
, DRO2, DRO3, DRO4, DRO5, DRO6, CAL, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16
, LINK17, LINK18, LINK19, LINK20, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input SPI1;
    input SPI2;
    input SPI3;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter inv_di_fclk1 = 1'b0;
    parameter inv_di_fclk2 = 1'b0;
    parameter latency1 = 1'b0;
    parameter latency2 = 1'b0;
    parameter location = "";
    parameter mode_cpath = "";
    parameter mode_epath = "";
    parameter mode_io_cal = 1'b0;
    parameter mode_rpath = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_tpath = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_CONTROL_U(ALCK1, ALCK2, ALCK3, LDSCK1, LDSCK2, LDSCK3, SWRX1CK, SWRX2CK, FCK1, FCK2, FDCK, CCK, DQ1CI1, DQ1CI2, DQ1CI3, DQ1CI4, DQ1CI5, DQ1CI6, DQ1CI7, DQ1CI8, DQ2CI1
, DQ2CI2, DQ2CI3, DQ2CI4, DQ2CI5, DQ2CI6, DQ2CI7, DQ2CI8, DQ3CI1, DQ3CI2, DQ3CI3, DQ3CI4, DQ3CI5, DQ3CI6, DQ3CI7, DQ3CI8, DQS1CI1, DQS1CI2, DQS1CI3, DQS1CI4, DQS1CI5, DQS1CI6
, DQS1CI7, DQS1CI8, DQS2CI1, DQS2CI2, DQS2CI3, DQS2CI4, DQS2CI5, DQS2CI6, DQS2CI7, DQS2CI8, DQS3CI1, DQS3CI2, DQS3CI3, DQS3CI4, DQS3CI5, DQS3CI6, DQS3CI7, DQS3CI8, LD1RN, LD2RN, LD3RN
, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DCRN, LE, SE, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3, DRA4, DRO1CSN
, DRO2CSN, DRO3CSN, DRI1CSN, DRI2CSN, DRI3CSN, DRDPA1CSN, DRDPA2CSN, DRDPA3CSN, DRCCSN, DRWDS, DRWEN, DRE, CA1P1, CA1P2, CA1P3, CA1P4, CA2P1, CA2P2, CA2P3, CA2P4, CA1N1
, CA1N2, CA1N3, CA1N4, CA2N1, CA2N2, CA2N3, CA2N4, CA1T1, CA1T2, CA1T3, CA1T4, CA2T1, CA2T2, CA2T3, CA2T4, CA1D1, CA1D2, CA1D3, CA1D4, CA1D5, CA1D6
, CA2D1, CA2D2, CA2D3, CA2D4, CA2D5, CA2D6, CKO1, CKO2, FLD, FLG, AL1D, AL2D, AL3D, AL1T, AL2T, AL3T, DCL, DRO1, DRO2, DRO3, DRO4
, DRO5, DRO6, LINK2, LINK3, LINK4, LINK5, LINK6, LINK7, LINK8, LINK9, LINK10, LINK11, LINK12, LINK13, LINK14, LINK15, LINK16, LINK17, LINK18, LINK19, LINK20
, LINK21, LINK22, LINK23, LINK24, LINK25, LINK26, LINK27, LINK28, LINK29, LINK30, LINK31, LINK32, LINK33, LINK34, LINK1);
    output AL1D;
    output AL1T;
    output AL2D;
    output AL2T;
    output AL3D;
    output AL3T;
    input ALCK1;
    input ALCK2;
    input ALCK3;
    input CA1D1;
    input CA1D2;
    input CA1D3;
    input CA1D4;
    input CA1D5;
    input CA1D6;
    input CA1N1;
    input CA1N2;
    input CA1N3;
    input CA1N4;
    input CA1P1;
    input CA1P2;
    input CA1P3;
    input CA1P4;
    input CA1T1;
    input CA1T2;
    input CA1T3;
    input CA1T4;
    input CA2D1;
    input CA2D2;
    input CA2D3;
    input CA2D4;
    input CA2D5;
    input CA2D6;
    input CA2N1;
    input CA2N2;
    input CA2N3;
    input CA2N4;
    input CA2P1;
    input CA2P2;
    input CA2P3;
    input CA2P4;
    input CA2T1;
    input CA2T2;
    input CA2T3;
    input CA2T4;
    input CCK;
    output CKO1;
    output CKO2;
    output DCL;
    input DCRN;
    input DQ1CI1;
    input DQ1CI2;
    input DQ1CI3;
    input DQ1CI4;
    input DQ1CI5;
    input DQ1CI6;
    input DQ1CI7;
    input DQ1CI8;
    input DQ2CI1;
    input DQ2CI2;
    input DQ2CI3;
    input DQ2CI4;
    input DQ2CI5;
    input DQ2CI6;
    input DQ2CI7;
    input DQ2CI8;
    input DQ3CI1;
    input DQ3CI2;
    input DQ3CI3;
    input DQ3CI4;
    input DQ3CI5;
    input DQ3CI6;
    input DQ3CI7;
    input DQ3CI8;
    input DQS1CI1;
    input DQS1CI2;
    input DQS1CI3;
    input DQS1CI4;
    input DQS1CI5;
    input DQS1CI6;
    input DQS1CI7;
    input DQS1CI8;
    input DQS2CI1;
    input DQS2CI2;
    input DQS2CI3;
    input DQS2CI4;
    input DQS2CI5;
    input DQS2CI6;
    input DQS2CI7;
    input DQS2CI8;
    input DQS3CI1;
    input DQS3CI2;
    input DQS3CI3;
    input DQS3CI4;
    input DQS3CI5;
    input DQS3CI6;
    input DQS3CI7;
    input DQS3CI8;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRCCSN;
    input DRDPA1CSN;
    input DRDPA2CSN;
    input DRDPA3CSN;
    input DRE;
    input DRI1;
    input DRI1CSN;
    input DRI2;
    input DRI2CSN;
    input DRI3;
    input DRI3CSN;
    input DRI4;
    input DRI5;
    input DRI6;
    output DRO1;
    input DRO1CSN;
    output DRO2;
    input DRO2CSN;
    output DRO3;
    input DRO3CSN;
    output DRO4;
    output DRO5;
    output DRO6;
    input DRWDS;
    input DRWEN;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    input FCK1;
    input FCK2;
    input FDCK;
    output FLD;
    output FLG;
    input FZ;
    input LD1RN;
    input LD2RN;
    input LD3RN;
    input LDSCK1;
    input LDSCK2;
    input LDSCK3;
    input LE;
    inout [41:0] LINK1;
    inout [41:0] LINK10;
    inout [41:0] LINK11;
    inout [41:0] LINK12;
    inout [41:0] LINK13;
    inout [41:0] LINK14;
    inout [41:0] LINK15;
    inout [41:0] LINK16;
    inout [41:0] LINK17;
    inout [41:0] LINK18;
    inout [41:0] LINK19;
    inout [41:0] LINK2;
    inout [41:0] LINK20;
    inout [41:0] LINK21;
    inout [41:0] LINK22;
    inout [41:0] LINK23;
    inout [41:0] LINK24;
    inout [41:0] LINK25;
    inout [41:0] LINK26;
    inout [41:0] LINK27;
    inout [41:0] LINK28;
    inout [41:0] LINK29;
    inout [41:0] LINK3;
    inout [41:0] LINK30;
    inout [41:0] LINK31;
    inout [41:0] LINK32;
    inout [41:0] LINK33;
    inout [41:0] LINK34;
    inout [41:0] LINK4;
    inout [41:0] LINK5;
    inout [41:0] LINK6;
    inout [41:0] LINK7;
    inout [41:0] LINK8;
    inout [41:0] LINK9;
    input SE;
    input SWRX1CK;
    input SWRX2CK;
    parameter cal_delay1 = "";
    parameter cal_delay2 = "";
    parameter div1 = 3'b000;
    parameter div2 = 3'b000;
    parameter div3 = 3'b000;
    parameter div_swrx1 = 3'b000;
    parameter div_swrx2 = 3'b000;
    parameter inv_ld_sck1 = 1'b0;
    parameter inv_ld_sck2 = 1'b0;
    parameter inv_ld_sck3 = 1'b0;
    parameter link_ld_12 = 1'b0;
    parameter link_ld_23 = 1'b0;
    parameter location = "";
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_side3 = 0;
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_dc_clk = 2'b00;
    parameter sel_ld_fck1 = 2'b00;
    parameter sel_ld_fck2 = 2'b00;
    parameter sel_ld_fck3 = 2'b00;
    parameter sel_sw_fck1 = 2'b00;
    parameter sel_sw_fck2 = 2'b00;
    parameter use_dc = 1'b0;
endmodule

(* blackbox *)
module NX_IOM_DRIVER(EI1, EI2, EI3, EI4, EI5, EL, ER, CI1, CI2, CI3, CI4, CI5, CL, CR, CTI, RI, RL, RR, CO, EO, RO1
, RO2, RO3, RO4, RO5, CTO, LINK);
    input CI1;
    input CI2;
    input CI3;
    input CI4;
    input CI5;
    input CL;
    output CO;
    input CR;
    input CTI;
    output CTO;
    input EI1;
    input EI2;
    input EI3;
    input EI4;
    input EI5;
    input EL;
    output EO;
    input ER;
    inout [41:0] LINK;
    input RI;
    input RL;
    output RO1;
    output RO2;
    output RO3;
    output RO4;
    output RO5;
    input RR;
    parameter chained = 1'b0;
    parameter cpath_edge = 1'b0;
    parameter cpath_init = 1'b0;
    parameter cpath_inv = 1'b0;
    parameter cpath_load = 1'b0;
    parameter cpath_mode = 4'b0000;
    parameter cpath_sync = 1'b0;
    parameter epath_dynamic = 1'b0;
    parameter epath_edge = 1'b0;
    parameter epath_init = 1'b0;
    parameter epath_load = 1'b0;
    parameter epath_mode = 4'b0000;
    parameter epath_sync = 1'b0;
    parameter location = "";
    parameter rpath_dynamic = 1'b0;
    parameter rpath_edge = 1'b0;
    parameter rpath_init = 1'b0;
    parameter rpath_load = 1'b0;
    parameter rpath_mode = 4'b0000;
    parameter rpath_sync = 1'b0;
    parameter symbol = "";
    parameter tpath_mode = 2'b00;
    parameter variant = "";
endmodule

(* blackbox *)
module NX_IOM_DRIVER_M(EI1, EI2, EI3, EI4, EI5, EL, ER, CI1, CI2, CI3, CI4, CI5, CL, CR, CTI, RI, RL, RR, CO, EO, RO1
, RO2, RO3, RO4, RO5, CTO, LINK);
    input CI1;
    input CI2;
    input CI3;
    input CI4;
    input CI5;
    input CL;
    output CO;
    input CR;
    input CTI;
    output CTO;
    input EI1;
    input EI2;
    input EI3;
    input EI4;
    input EI5;
    input EL;
    output EO;
    input ER;
    inout [41:0] LINK;
    input RI;
    input RL;
    output RO1;
    output RO2;
    output RO3;
    output RO4;
    output RO5;
    input RR;
    parameter chained = 1'b0;
    parameter cpath_edge = 1'b0;
    parameter cpath_init = 1'b0;
    parameter cpath_inv = 1'b0;
    parameter cpath_load = 1'b0;
    parameter cpath_mode = 4'b0000;
    parameter cpath_sync = 1'b0;
    parameter epath_dynamic = 1'b0;
    parameter epath_edge = 1'b0;
    parameter epath_init = 1'b0;
    parameter epath_load = 1'b0;
    parameter epath_mode = 4'b0000;
    parameter epath_sync = 1'b0;
    parameter location = "";
    parameter rpath_dynamic = 1'b0;
    parameter rpath_edge = 1'b0;
    parameter rpath_init = 1'b0;
    parameter rpath_load = 1'b0;
    parameter rpath_mode = 4'b0000;
    parameter rpath_sync = 1'b0;
    parameter symbol = "";
    parameter tpath_mode = 2'b00;
    parameter variant = "";
endmodule

(* blackbox *)
module NX_IOM_DRIVER_U(EI1, EI2, EI3, EI4, EI5, EI6, EI7, EI8, EL, ER, CI1, CL, CR, RI, RL, RR, CO, CTI, CTO, EO, RO1
, RO2, RO3, RO4, RO5, RO6, RO7, RO8, LINK);
    input CI1;
    input CL;
    output CO;
    input CR;
    input CTI;
    output CTO;
    input EI1;
    input EI2;
    input EI3;
    input EI4;
    input EI5;
    input EI6;
    input EI7;
    input EI8;
    input EL;
    output EO;
    input ER;
    inout [41:0] LINK;
    input RI;
    input RL;
    output RO1;
    output RO2;
    output RO3;
    output RO4;
    output RO5;
    output RO6;
    output RO7;
    output RO8;
    input RR;
    parameter chained = 1'b0;
    parameter cpath_edge = 1'b0;
    parameter cpath_init = 1'b0;
    parameter cpath_inv = 1'b0;
    parameter cpath_load = 1'b0;
    parameter cpath_mode = 4'b0000;
    parameter cpath_sync = 1'b0;
    parameter cpath_type = 1'b0;
    parameter epath_dynamic = 1'b0;
    parameter epath_edge = 1'b0;
    parameter epath_init = 1'b0;
    parameter epath_load = 1'b0;
    parameter epath_mode = 4'b0000;
    parameter epath_sync = 1'b0;
    parameter epath_type = 1'b0;
    parameter location = "";
    parameter rpath_dynamic = 1'b0;
    parameter rpath_edge = 1'b0;
    parameter rpath_init = 1'b0;
    parameter rpath_load = 1'b0;
    parameter rpath_mode = 4'b0000;
    parameter rpath_sync = 1'b0;
    parameter rpath_type = 1'b0;
    parameter symbol = "";
    parameter tpath_mode = 1'b0;
endmodule

(* blackbox *)
module NX_IOM_L(RTCK1, RRCK1, WTCK1, WRCK1, RTCK2, RRCK2, WTCK2, WRCK2, CTCK, CCK, DCK, C1TW, C1TS, C1RW1, C1RW2, C1RW3, C1RNE, C1RS, C2TW, C2TS, C2RW1
, C2RW2, C2RW3, C2RNE, C2RS, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DC, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3
, DRA4, DRA5, DRA6, DRL, DOS, DOG, DIS, DIG, DPAS, DPAG, DQSS, DQSG, DS1, DS2, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CAP1
, CAP2, CAP3, CAP4, CAN1, CAN2, CAN3, CAN4, CAT1, CAT2, CAT3, CAT4, CKO1, CKO2, FLD, FLG, C1RED, C2RED, DRO1, DRO2, DRO3, DRO4
, DRO5, DRO6, CAL, P1CI1, P1CL, P1CR, P1CO, P1CTI, P1CTO, P1EI1, P1EI2, P1EI3, P1EI4, P1EI5, P1EL, P1ER, P1EO, P1RI, P1RL, P1RR, P1RO1
, P1RO2, P1RO3, P1RO4, P1RO5, P2CI1, P2CL, P2CR, P2CO, P2CTI, P2CTO, P2EI1, P2EI2, P2EI3, P2EI4, P2EI5, P2EL, P2ER, P2EO, P2RI, P2RL, P2RR
, P2RO1, P2RO2, P2RO3, P2RO4, P2RO5, P3CI1, P3CL, P3CR, P3CO, P3CTI, P3CTO, P3EI1, P3EI2, P3EI3, P3EI4, P3EI5, P3EL, P3ER, P3EO, P3RI, P3RL
, P3RR, P3RO1, P3RO2, P3RO3, P3RO4, P3RO5, P4CI1, P4CL, P4CR, P4CO, P4CTI, P4CTO, P4EI1, P4EI2, P4EI3, P4EI4, P4EI5, P4EL, P4ER, P4EO, P4RI
, P4RL, P4RR, P4RO1, P4RO2, P4RO3, P4RO4, P4RO5, P5CI1, P5CI2, P5CI3, P5CI4, P5CI5, P5CL, P5CR, P5CO, P5CTI, P5CTO, P5EI1, P5EI2, P5EI3, P5EI4
, P5EI5, P5EL, P5ER, P5EO, P5RI, P5RL, P5RR, P5RO1, P5RO2, P5RO3, P5RO4, P5RO5, P6CI1, P6CL, P6CR, P6CO, P6CTI, P6CTO, P6EI1, P6EI2, P6EI3
, P6EI4, P6EI5, P6EL, P6ER, P6EO, P6RI, P6RL, P6RR, P6RO1, P6RO2, P6RO3, P6RO4, P6RO5, P7CI1, P7CL, P7CR, P7CO, P7CTI, P7CTO, P7EI1, P7EI2
, P7EI3, P7EI4, P7EI5, P7EL, P7ER, P7EO, P7RI, P7RL, P7RR, P7RO1, P7RO2, P7RO3, P7RO4, P7RO5, P8CI1, P8CL, P8CR, P8CO, P8CTI, P8CTO, P8EI1
, P8EI2, P8EI3, P8EI4, P8EI5, P8EL, P8ER, P8EO, P8RI, P8RL, P8RR, P8RO1, P8RO2, P8RO3, P8RO4, P8RO5, P9CI1, P9CL, P9CR, P9CO, P9CTI, P9CTO
, P9EI1, P9EI2, P9EI3, P9EI4, P9EI5, P9EL, P9ER, P9EO, P9RI, P9RL, P9RR, P9RO1, P9RO2, P9RO3, P9RO4, P9RO5, P10CI1, P10CL, P10CR, P10CO, P10CTI
, P10CTO, P10EI1, P10EI2, P10EI3, P10EI4, P10EI5, P10EL, P10ER, P10EO, P10RI, P10RL, P10RR, P10RO1, P10RO2, P10RO3, P10RO4, P10RO5, P11CI1, P11CL, P11CR, P11CO
, P11CTI, P11CTO, P11EI1, P11EI2, P11EI3, P11EI4, P11EI5, P11EL, P11ER, P11EO, P11RI, P11RL, P11RR, P11RO1, P11RO2, P11RO3, P11RO4, P11RO5, P12CI1, P12CL, P12CR
, P12CO, P12CTI, P12CTO, P12EI1, P12EI2, P12EI3, P12EI4, P12EI5, P12EL, P12ER, P12EO, P12RI, P12RL, P12RR, P12RO1, P12RO2, P12RO3, P12RO4, P12RO5, P13CI1, P13CL
, P13CR, P13CO, P13CTI, P13CTO, P13EI1, P13EI2, P13EI3, P13EI4, P13EI5, P13EL, P13ER, P13EO, P13RI, P13RL, P13RR, P13RO1, P13RO2, P13RO3, P13RO4, P13RO5, P14CI1
, P14CL, P14CR, P14CO, P14CTI, P14CTO, P14EI1, P14EI2, P14EI3, P14EI4, P14EI5, P14EL, P14ER, P14EO, P14RI, P14RL, P14RR, P14RO1, P14RO2, P14RO3, P14RO4, P14RO5
, P15CI1, P15CL, P15CR, P15CO, P15CTI, P15CTO, P15EI1, P15EI2, P15EI3, P15EI4, P15EI5, P15EL, P15ER, P15EO, P15RI, P15RL, P15RR, P15RO1, P15RO2, P15RO3, P15RO4
, P15RO5, P16CI1, P16CL, P16CR, P16CO, P16CTI, P16CTO, P16EI1, P16EI2, P16EI3, P16EI4, P16EI5, P16EL, P16ER, P16EO, P16RI, P16RL, P16RR, P16RO1, P16RO2, P16RO3
, P16RO4, P16RO5, P17CI1, P17CL, P17CR, P17CO, P17CTI, P17CTO, P17EI1, P17EI2, P17EI3, P17EI4, P17EI5, P17EL, P17ER, P17EO, P17RI, P17RL, P17RR, P17RO1, P17RO2
, P17RO3, P17RO4, P17RO5, P18CI1, P18CL, P18CR, P18CO, P18CTI, P18CTO, P18EI1, P18EI2, P18EI3, P18EI4, P18EI5, P18EL, P18ER, P18EO, P18RI, P18RL, P18RR, P18RO1
, P18RO2, P18RO3, P18RO4, P18RO5, P19CI1, P19CL, P19CR, P19CO, P19CTI, P19CTO, P19EI1, P19EI2, P19EI3, P19EI4, P19EI5, P19EL, P19ER, P19EO, P19RI, P19RL, P19RR
, P19RO1, P19RO2, P19RO3, P19RO4, P19RO5, P20CI1, P20CL, P20CR, P20CO, P20CTI, P20CTO, P20EI1, P20EI2, P20EI3, P20EI4, P20EI5, P20EL, P20ER, P20EO, P20RI, P20RL
, P20RR, P20RO1, P20RO2, P20RO3, P20RO4, P20RO5, P21CI1, P21CL, P21CR, P21CO, P21CTI, P21CTO, P21EI1, P21EI2, P21EI3, P21EI4, P21EI5, P21EL, P21ER, P21EO, P21RI
, P21RL, P21RR, P21RO1, P21RO2, P21RO3, P21RO4, P21RO5, P22CI1, P22CL, P22CR, P22CO, P22CTI, P22CTO, P22EI1, P22EI2, P22EI3, P22EI4, P22EI5, P22EL, P22ER, P22EO
, P22RI, P22RL, P22RR, P22RO1, P22RO2, P22RO3, P22RO4, P22RO5, P23CI1, P23CL, P23CR, P23CO, P23CTI, P23CTO, P23EI1, P23EI2, P23EI3, P23EI4, P23EI5, P23EL, P23ER
, P23EO, P23RI, P23RL, P23RR, P23RO1, P23RO2, P23RO3, P23RO4, P23RO5, P24CI1, P24CL, P24CR, P24CO, P24CTI, P24CTO, P24EI1, P24EI2, P24EI3, P24EI4, P24EI5, P24EL
, P24ER, P24EO, P24RI, P24RL, P24RR, P24RO1, P24RO2, P24RO3, P24RO4, P24RO5, P25CI1, P25CL, P25CR, P25CO, P25CTI, P25CTO, P25EI1, P25EI2, P25EI3, P25EI4, P25EI5
, P25EL, P25ER, P25EO, P25RI, P25RL, P25RR, P25RO1, P25RO2, P25RO3, P25RO4, P25RO5, P26CI1, P26CL, P26CR, P26CO, P26CTI, P26CTO, P26EI1, P26EI2, P26EI3, P26EI4
, P26EI5, P26EL, P26ER, P26EO, P26RI, P26RL, P26RR, P26RO1, P26RO2, P26RO3, P26RO4, P26RO5, P27CI1, P27CL, P27CR, P27CO, P27CTI, P27CTO, P27EI1, P27EI2, P27EI3
, P27EI4, P27EI5, P27EL, P27ER, P27EO, P27RI, P27RL, P27RR, P27RO1, P27RO2, P27RO3, P27RO4, P27RO5, P28CI1, P28CL, P28CR, P28CO, P28CTI, P28CTO, P28EI1, P28EI2
, P28EI3, P28EI4, P28EI5, P28EL, P28ER, P28EO, P28RI, P28RL, P28RR, P28RO1, P28RO2, P28RO3, P28RO4, P28RO5, P29CI1, P29CI2, P29CI3, P29CI4, P29CI5, P29CL, P29CR
, P29CO, P29CTI, P29CTO, P29EI1, P29EI2, P29EI3, P29EI4, P29EI5, P29EL, P29ER, P29EO, P29RI, P29RL, P29RR, P29RO1, P29RO2, P29RO3, P29RO4, P29RO5, P30CI1, P30CL
, P30CR, P30CO, P30CTI, P30CTO, P30EI1, P30EI2, P30EI3, P30EI4, P30EI5, P30EL, P30ER, P30EO, P30RI, P30RL, P30RR, P30RO1, P30RO2, P30RO3, P30RO4, P30RO5, P31CI1
, P31CL, P31CR, P31CO, P31CTI, P31CTO, P31EI1, P31EI2, P31EI3, P31EI4, P31EI5, P31EL, P31ER, P31EO, P31RI, P31RL, P31RR, P31RO1, P31RO2, P31RO3, P31RO4, P31RO5
, P32CI1, P32CL, P32CR, P32CO, P32CTI, P32CTO, P32EI1, P32EI2, P32EI3, P32EI4, P32EI5, P32EL, P32ER, P32EO, P32RI, P32RL, P32RR, P32RO1, P32RO2, P32RO3, P32RO4
, P32RO5, P33CI1, P33CL, P33CR, P33CO, P33CTI, P33CTO, P33EI1, P33EI2, P33EI3, P33EI4, P33EI5, P33EL, P33ER, P33EO, P33RI, P33RL, P33RR, P33RO1, P33RO2, P33RO3
, P33RO4, P33RO5, P34CI1, P34CL, P34CR, P34CO, P34CTI, P34CTO, P34EI1, P34EI2, P34EI3, P34EI4, P34EI5, P34EL, P34ER, P34EO, P34RI, P34RL, P34RR, P34RO1, P34RO2
, P34RO3, P34RO4, P34RO5);
    output C1RED;
    input C1RNE;
    input C1RS;
    input C1RW1;
    input C1RW2;
    input C1RW3;
    input C1TS;
    input C1TW;
    output C2RED;
    input C2RNE;
    input C2RS;
    input C2RW1;
    input C2RW2;
    input C2RW3;
    input C2TS;
    input C2TW;
    input CAD1;
    input CAD2;
    input CAD3;
    input CAD4;
    input CAD5;
    input CAD6;
    output CAL;
    input CAN1;
    input CAN2;
    input CAN3;
    input CAN4;
    input CAP1;
    input CAP2;
    input CAP3;
    input CAP4;
    input CAT1;
    input CAT2;
    input CAT3;
    input CAT4;
    input CCK;
    output CKO1;
    output CKO2;
    input CTCK;
    input DC;
    input DCK;
    input DIG;
    input DIS;
    input DOG;
    input DOS;
    input DPAG;
    input DPAS;
    input DQSG;
    input DQSS;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRA5;
    input DRA6;
    input DRI1;
    input DRI2;
    input DRI3;
    input DRI4;
    input DRI5;
    input DRI6;
    input DRL;
    output DRO1;
    output DRO2;
    output DRO3;
    output DRO4;
    output DRO5;
    output DRO6;
    input DS1;
    input DS2;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    output FLD;
    output FLG;
    input FZ;
    input P10CI1;
    input P10CL;
    output P10CO;
    input P10CR;
    input P10CTI;
    output P10CTO;
    input P10EI1;
    input P10EI2;
    input P10EI3;
    input P10EI4;
    input P10EI5;
    input P10EL;
    output P10EO;
    input P10ER;
    input P10RI;
    input P10RL;
    output P10RO1;
    output P10RO2;
    output P10RO3;
    output P10RO4;
    output P10RO5;
    input P10RR;
    input P11CI1;
    input P11CL;
    output P11CO;
    input P11CR;
    input P11CTI;
    output P11CTO;
    input P11EI1;
    input P11EI2;
    input P11EI3;
    input P11EI4;
    input P11EI5;
    input P11EL;
    output P11EO;
    input P11ER;
    input P11RI;
    input P11RL;
    output P11RO1;
    output P11RO2;
    output P11RO3;
    output P11RO4;
    output P11RO5;
    input P11RR;
    input P12CI1;
    input P12CL;
    output P12CO;
    input P12CR;
    input P12CTI;
    output P12CTO;
    input P12EI1;
    input P12EI2;
    input P12EI3;
    input P12EI4;
    input P12EI5;
    input P12EL;
    output P12EO;
    input P12ER;
    input P12RI;
    input P12RL;
    output P12RO1;
    output P12RO2;
    output P12RO3;
    output P12RO4;
    output P12RO5;
    input P12RR;
    input P13CI1;
    input P13CL;
    output P13CO;
    input P13CR;
    input P13CTI;
    output P13CTO;
    input P13EI1;
    input P13EI2;
    input P13EI3;
    input P13EI4;
    input P13EI5;
    input P13EL;
    output P13EO;
    input P13ER;
    input P13RI;
    input P13RL;
    output P13RO1;
    output P13RO2;
    output P13RO3;
    output P13RO4;
    output P13RO5;
    input P13RR;
    input P14CI1;
    input P14CL;
    output P14CO;
    input P14CR;
    input P14CTI;
    output P14CTO;
    input P14EI1;
    input P14EI2;
    input P14EI3;
    input P14EI4;
    input P14EI5;
    input P14EL;
    output P14EO;
    input P14ER;
    input P14RI;
    input P14RL;
    output P14RO1;
    output P14RO2;
    output P14RO3;
    output P14RO4;
    output P14RO5;
    input P14RR;
    input P15CI1;
    input P15CL;
    output P15CO;
    input P15CR;
    input P15CTI;
    output P15CTO;
    input P15EI1;
    input P15EI2;
    input P15EI3;
    input P15EI4;
    input P15EI5;
    input P15EL;
    output P15EO;
    input P15ER;
    input P15RI;
    input P15RL;
    output P15RO1;
    output P15RO2;
    output P15RO3;
    output P15RO4;
    output P15RO5;
    input P15RR;
    input P16CI1;
    input P16CL;
    output P16CO;
    input P16CR;
    input P16CTI;
    output P16CTO;
    input P16EI1;
    input P16EI2;
    input P16EI3;
    input P16EI4;
    input P16EI5;
    input P16EL;
    output P16EO;
    input P16ER;
    input P16RI;
    input P16RL;
    output P16RO1;
    output P16RO2;
    output P16RO3;
    output P16RO4;
    output P16RO5;
    input P16RR;
    input P17CI1;
    input P17CL;
    output P17CO;
    input P17CR;
    input P17CTI;
    output P17CTO;
    input P17EI1;
    input P17EI2;
    input P17EI3;
    input P17EI4;
    input P17EI5;
    input P17EL;
    output P17EO;
    input P17ER;
    input P17RI;
    input P17RL;
    output P17RO1;
    output P17RO2;
    output P17RO3;
    output P17RO4;
    output P17RO5;
    input P17RR;
    input P18CI1;
    input P18CL;
    output P18CO;
    input P18CR;
    input P18CTI;
    output P18CTO;
    input P18EI1;
    input P18EI2;
    input P18EI3;
    input P18EI4;
    input P18EI5;
    input P18EL;
    output P18EO;
    input P18ER;
    input P18RI;
    input P18RL;
    output P18RO1;
    output P18RO2;
    output P18RO3;
    output P18RO4;
    output P18RO5;
    input P18RR;
    input P19CI1;
    input P19CL;
    output P19CO;
    input P19CR;
    input P19CTI;
    output P19CTO;
    input P19EI1;
    input P19EI2;
    input P19EI3;
    input P19EI4;
    input P19EI5;
    input P19EL;
    output P19EO;
    input P19ER;
    input P19RI;
    input P19RL;
    output P19RO1;
    output P19RO2;
    output P19RO3;
    output P19RO4;
    output P19RO5;
    input P19RR;
    input P1CI1;
    input P1CL;
    output P1CO;
    input P1CR;
    input P1CTI;
    output P1CTO;
    input P1EI1;
    input P1EI2;
    input P1EI3;
    input P1EI4;
    input P1EI5;
    input P1EL;
    output P1EO;
    input P1ER;
    input P1RI;
    input P1RL;
    output P1RO1;
    output P1RO2;
    output P1RO3;
    output P1RO4;
    output P1RO5;
    input P1RR;
    input P20CI1;
    input P20CL;
    output P20CO;
    input P20CR;
    input P20CTI;
    output P20CTO;
    input P20EI1;
    input P20EI2;
    input P20EI3;
    input P20EI4;
    input P20EI5;
    input P20EL;
    output P20EO;
    input P20ER;
    input P20RI;
    input P20RL;
    output P20RO1;
    output P20RO2;
    output P20RO3;
    output P20RO4;
    output P20RO5;
    input P20RR;
    input P21CI1;
    input P21CL;
    output P21CO;
    input P21CR;
    input P21CTI;
    output P21CTO;
    input P21EI1;
    input P21EI2;
    input P21EI3;
    input P21EI4;
    input P21EI5;
    input P21EL;
    output P21EO;
    input P21ER;
    input P21RI;
    input P21RL;
    output P21RO1;
    output P21RO2;
    output P21RO3;
    output P21RO4;
    output P21RO5;
    input P21RR;
    input P22CI1;
    input P22CL;
    output P22CO;
    input P22CR;
    input P22CTI;
    output P22CTO;
    input P22EI1;
    input P22EI2;
    input P22EI3;
    input P22EI4;
    input P22EI5;
    input P22EL;
    output P22EO;
    input P22ER;
    input P22RI;
    input P22RL;
    output P22RO1;
    output P22RO2;
    output P22RO3;
    output P22RO4;
    output P22RO5;
    input P22RR;
    input P23CI1;
    input P23CL;
    output P23CO;
    input P23CR;
    input P23CTI;
    output P23CTO;
    input P23EI1;
    input P23EI2;
    input P23EI3;
    input P23EI4;
    input P23EI5;
    input P23EL;
    output P23EO;
    input P23ER;
    input P23RI;
    input P23RL;
    output P23RO1;
    output P23RO2;
    output P23RO3;
    output P23RO4;
    output P23RO5;
    input P23RR;
    input P24CI1;
    input P24CL;
    output P24CO;
    input P24CR;
    input P24CTI;
    output P24CTO;
    input P24EI1;
    input P24EI2;
    input P24EI3;
    input P24EI4;
    input P24EI5;
    input P24EL;
    output P24EO;
    input P24ER;
    input P24RI;
    input P24RL;
    output P24RO1;
    output P24RO2;
    output P24RO3;
    output P24RO4;
    output P24RO5;
    input P24RR;
    input P25CI1;
    input P25CL;
    output P25CO;
    input P25CR;
    input P25CTI;
    output P25CTO;
    input P25EI1;
    input P25EI2;
    input P25EI3;
    input P25EI4;
    input P25EI5;
    input P25EL;
    output P25EO;
    input P25ER;
    input P25RI;
    input P25RL;
    output P25RO1;
    output P25RO2;
    output P25RO3;
    output P25RO4;
    output P25RO5;
    input P25RR;
    input P26CI1;
    input P26CL;
    output P26CO;
    input P26CR;
    input P26CTI;
    output P26CTO;
    input P26EI1;
    input P26EI2;
    input P26EI3;
    input P26EI4;
    input P26EI5;
    input P26EL;
    output P26EO;
    input P26ER;
    input P26RI;
    input P26RL;
    output P26RO1;
    output P26RO2;
    output P26RO3;
    output P26RO4;
    output P26RO5;
    input P26RR;
    input P27CI1;
    input P27CL;
    output P27CO;
    input P27CR;
    input P27CTI;
    output P27CTO;
    input P27EI1;
    input P27EI2;
    input P27EI3;
    input P27EI4;
    input P27EI5;
    input P27EL;
    output P27EO;
    input P27ER;
    input P27RI;
    input P27RL;
    output P27RO1;
    output P27RO2;
    output P27RO3;
    output P27RO4;
    output P27RO5;
    input P27RR;
    input P28CI1;
    input P28CL;
    output P28CO;
    input P28CR;
    input P28CTI;
    output P28CTO;
    input P28EI1;
    input P28EI2;
    input P28EI3;
    input P28EI4;
    input P28EI5;
    input P28EL;
    output P28EO;
    input P28ER;
    input P28RI;
    input P28RL;
    output P28RO1;
    output P28RO2;
    output P28RO3;
    output P28RO4;
    output P28RO5;
    input P28RR;
    input P29CI1;
    input P29CI2;
    input P29CI3;
    input P29CI4;
    input P29CI5;
    input P29CL;
    output P29CO;
    input P29CR;
    input P29CTI;
    output P29CTO;
    input P29EI1;
    input P29EI2;
    input P29EI3;
    input P29EI4;
    input P29EI5;
    input P29EL;
    output P29EO;
    input P29ER;
    input P29RI;
    input P29RL;
    output P29RO1;
    output P29RO2;
    output P29RO3;
    output P29RO4;
    output P29RO5;
    input P29RR;
    input P2CI1;
    input P2CL;
    output P2CO;
    input P2CR;
    input P2CTI;
    output P2CTO;
    input P2EI1;
    input P2EI2;
    input P2EI3;
    input P2EI4;
    input P2EI5;
    input P2EL;
    output P2EO;
    input P2ER;
    input P2RI;
    input P2RL;
    output P2RO1;
    output P2RO2;
    output P2RO3;
    output P2RO4;
    output P2RO5;
    input P2RR;
    input P30CI1;
    input P30CL;
    output P30CO;
    input P30CR;
    input P30CTI;
    output P30CTO;
    input P30EI1;
    input P30EI2;
    input P30EI3;
    input P30EI4;
    input P30EI5;
    input P30EL;
    output P30EO;
    input P30ER;
    input P30RI;
    input P30RL;
    output P30RO1;
    output P30RO2;
    output P30RO3;
    output P30RO4;
    output P30RO5;
    input P30RR;
    input P31CI1;
    input P31CL;
    output P31CO;
    input P31CR;
    input P31CTI;
    output P31CTO;
    input P31EI1;
    input P31EI2;
    input P31EI3;
    input P31EI4;
    input P31EI5;
    input P31EL;
    output P31EO;
    input P31ER;
    input P31RI;
    input P31RL;
    output P31RO1;
    output P31RO2;
    output P31RO3;
    output P31RO4;
    output P31RO5;
    input P31RR;
    input P32CI1;
    input P32CL;
    output P32CO;
    input P32CR;
    input P32CTI;
    output P32CTO;
    input P32EI1;
    input P32EI2;
    input P32EI3;
    input P32EI4;
    input P32EI5;
    input P32EL;
    output P32EO;
    input P32ER;
    input P32RI;
    input P32RL;
    output P32RO1;
    output P32RO2;
    output P32RO3;
    output P32RO4;
    output P32RO5;
    input P32RR;
    input P33CI1;
    input P33CL;
    output P33CO;
    input P33CR;
    input P33CTI;
    output P33CTO;
    input P33EI1;
    input P33EI2;
    input P33EI3;
    input P33EI4;
    input P33EI5;
    input P33EL;
    output P33EO;
    input P33ER;
    input P33RI;
    input P33RL;
    output P33RO1;
    output P33RO2;
    output P33RO3;
    output P33RO4;
    output P33RO5;
    input P33RR;
    input P34CI1;
    input P34CL;
    output P34CO;
    input P34CR;
    input P34CTI;
    output P34CTO;
    input P34EI1;
    input P34EI2;
    input P34EI3;
    input P34EI4;
    input P34EI5;
    input P34EL;
    output P34EO;
    input P34ER;
    input P34RI;
    input P34RL;
    output P34RO1;
    output P34RO2;
    output P34RO3;
    output P34RO4;
    output P34RO5;
    input P34RR;
    input P3CI1;
    input P3CL;
    output P3CO;
    input P3CR;
    input P3CTI;
    output P3CTO;
    input P3EI1;
    input P3EI2;
    input P3EI3;
    input P3EI4;
    input P3EI5;
    input P3EL;
    output P3EO;
    input P3ER;
    input P3RI;
    input P3RL;
    output P3RO1;
    output P3RO2;
    output P3RO3;
    output P3RO4;
    output P3RO5;
    input P3RR;
    input P4CI1;
    input P4CL;
    output P4CO;
    input P4CR;
    input P4CTI;
    output P4CTO;
    input P4EI1;
    input P4EI2;
    input P4EI3;
    input P4EI4;
    input P4EI5;
    input P4EL;
    output P4EO;
    input P4ER;
    input P4RI;
    input P4RL;
    output P4RO1;
    output P4RO2;
    output P4RO3;
    output P4RO4;
    output P4RO5;
    input P4RR;
    input P5CI1;
    input P5CI2;
    input P5CI3;
    input P5CI4;
    input P5CI5;
    input P5CL;
    output P5CO;
    input P5CR;
    input P5CTI;
    output P5CTO;
    input P5EI1;
    input P5EI2;
    input P5EI3;
    input P5EI4;
    input P5EI5;
    input P5EL;
    output P5EO;
    input P5ER;
    input P5RI;
    input P5RL;
    output P5RO1;
    output P5RO2;
    output P5RO3;
    output P5RO4;
    output P5RO5;
    input P5RR;
    input P6CI1;
    input P6CL;
    output P6CO;
    input P6CR;
    input P6CTI;
    output P6CTO;
    input P6EI1;
    input P6EI2;
    input P6EI3;
    input P6EI4;
    input P6EI5;
    input P6EL;
    output P6EO;
    input P6ER;
    input P6RI;
    input P6RL;
    output P6RO1;
    output P6RO2;
    output P6RO3;
    output P6RO4;
    output P6RO5;
    input P6RR;
    input P7CI1;
    input P7CL;
    output P7CO;
    input P7CR;
    input P7CTI;
    output P7CTO;
    input P7EI1;
    input P7EI2;
    input P7EI3;
    input P7EI4;
    input P7EI5;
    input P7EL;
    output P7EO;
    input P7ER;
    input P7RI;
    input P7RL;
    output P7RO1;
    output P7RO2;
    output P7RO3;
    output P7RO4;
    output P7RO5;
    input P7RR;
    input P8CI1;
    input P8CL;
    output P8CO;
    input P8CR;
    input P8CTI;
    output P8CTO;
    input P8EI1;
    input P8EI2;
    input P8EI3;
    input P8EI4;
    input P8EI5;
    input P8EL;
    output P8EO;
    input P8ER;
    input P8RI;
    input P8RL;
    output P8RO1;
    output P8RO2;
    output P8RO3;
    output P8RO4;
    output P8RO5;
    input P8RR;
    input P9CI1;
    input P9CL;
    output P9CO;
    input P9CR;
    input P9CTI;
    output P9CTO;
    input P9EI1;
    input P9EI2;
    input P9EI3;
    input P9EI4;
    input P9EI5;
    input P9EL;
    output P9EO;
    input P9ER;
    input P9RI;
    input P9RL;
    output P9RO1;
    output P9RO2;
    output P9RO3;
    output P9RO4;
    output P9RO5;
    input P9RR;
    input RRCK1;
    input RRCK2;
    input RTCK1;
    input RTCK2;
    input WRCK1;
    input WRCK2;
    input WTCK1;
    input WTCK2;
    parameter div_rx1 = 4'b0000;
    parameter div_rx2 = 4'b0000;
    parameter div_tx1 = 4'b0000;
    parameter div_tx2 = 4'b0000;
    parameter mode_io_cal = 1'b0;
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter pads_dict = "";
    parameter pads_path = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_clkr_rx1 = 1'b0;
    parameter sel_clkr_rx2 = 1'b0;
    parameter sel_clkw_rx1 = 2'b00;
    parameter sel_clkw_rx2 = 2'b00;
endmodule

(* blackbox *)
module NX_IOM_SERDES(RTCK, WRCK, WTCK, RRCK, TRST, RRST, CTCK, DCK, DRL, DIG, FZ, FLD, FLG, DS, DRA, DRI, DRO, DID, LINKN, LINKP);
    input CTCK;
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINKN;
    inout [41:0] LINKP;
    input RRCK;
    input RRST;
    input RTCK;
    input TRST;
    input WRCK;
    input WTCK;
    parameter data_size = 5;
    parameter location = "";
endmodule

(* blackbox *)
module NX_IOM_SERDES_M(RTCK, WRCK, WTCK, RRCK, TRST, RRST, CTCK, DCK, DRL, DIG, FZ, FLD, FLG, DS, DRA, DRI, DRO, DID, LINKN, LINKP);
    input CTCK;
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    output FLD;
    output FLG;
    input FZ;
    inout [41:0] LINKN;
    inout [41:0] LINKP;
    input RRCK;
    input RRST;
    input RTCK;
    input TRST;
    input WRCK;
    input WTCK;
    parameter data_size = 5;
    parameter location = "";
endmodule

(* blackbox *)
module NX_IOM_SERDES_U(FCK, SCK, LDRN, DRWDS, DRWEN, DRE, FZ, ALD, ALT, FLD, FLG, LINK, DRA, DRI, DRO, DID, DRIN, DRDN, FA, DRON);
    output ALD;
    output ALT;
    output [5:0] DID;
    input [3:0] DRA;
    input [2:0] DRDN;
    input DRE;
    input [5:0] DRI;
    input [2:0] DRIN;
    output [5:0] DRO;
    input [2:0] DRON;
    input DRWDS;
    input DRWEN;
    input [5:0] FA;
    input FCK;
    output FLD;
    output FLG;
    input FZ;
    input LDRN;
    inout [41:0] LINK;
    input SCK;
    parameter data_size = 5;
    parameter location = "";
endmodule

(* blackbox *)
module NX_IOM_U(ALCK1, ALCK2, ALCK3, LDSCK1, LDSCK2, LDSCK3, SWRX1CK, SWRX2CK, FCK1, FCK2, FDCK, CCK, DQ1CI1, DQ1CI2, DQ1CI3, DQ1CI4, DQ1CI5, DQ1CI6, DQ1CI7, DQ1CI8, DQ2CI1
, DQ2CI2, DQ2CI3, DQ2CI4, DQ2CI5, DQ2CI6, DQ2CI7, DQ2CI8, DQ3CI1, DQ3CI2, DQ3CI3, DQ3CI4, DQ3CI5, DQ3CI6, DQ3CI7, DQ3CI8, DQS1CI1, DQS1CI2, DQS1CI3, DQS1CI4, DQS1CI5, DQS1CI6
, DQS1CI7, DQS1CI8, DQS2CI1, DQS2CI2, DQS2CI3, DQS2CI4, DQS2CI5, DQS2CI6, DQS2CI7, DQS2CI8, DQS3CI1, DQS3CI2, DQS3CI3, DQS3CI4, DQS3CI5, DQS3CI6, DQS3CI7, DQS3CI8, LD1RN, LD2RN, LD3RN
, FA1, FA2, FA3, FA4, FA5, FA6, FZ, DCRN, LE, SE, DRI1, DRI2, DRI3, DRI4, DRI5, DRI6, DRA1, DRA2, DRA3, DRA4, DRO1CSN
, DRO2CSN, DRO3CSN, DRI1CSN, DRI2CSN, DRI3CSN, DRDPA1CSN, DRDPA2CSN, DRDPA3CSN, DRCCSN, DRWDS, DRWEN, DRE, CA1P1, CA1P2, CA1P3, CA1P4, CA2P1, CA2P2, CA2P3, CA2P4, CA1N1
, CA1N2, CA1N3, CA1N4, CA2N1, CA2N2, CA2N3, CA2N4, CA1T1, CA1T2, CA1T3, CA1T4, CA2T1, CA2T2, CA2T3, CA2T4, CA1D1, CA1D2, CA1D3, CA1D4, CA1D5, CA1D6
, CA2D1, CA2D2, CA2D3, CA2D4, CA2D5, CA2D6, CKO1, CKO2, FLD, FLG, AL1D, AL2D, AL3D, AL1T, AL2T, AL3T, DCL, DRO1, DRO2, DRO3, DRO4
, DRO5, DRO6, P1CI1, P1CL, P1CR, P1CO, P1CTI, P1CTO, P1EI1, P1EI2, P1EI3, P1EI4, P1EI5, P1EI6, P1EI7, P1EI8, P1EL, P1ER, P1EO, P1RI, P1RL
, P1RR, P1RO1, P1RO2, P1RO3, P1RO4, P1RO5, P1RO6, P1RO7, P1RO8, P2CI1, P2CL, P2CR, P2CO, P2CTI, P2CTO, P2EI1, P2EI2, P2EI3, P2EI4, P2EI5, P2EI6
, P2EI7, P2EI8, P2EL, P2ER, P2EO, P2RI, P2RL, P2RR, P2RO1, P2RO2, P2RO3, P2RO4, P2RO5, P2RO6, P2RO7, P2RO8, P3CI1, P3CL, P3CR, P3CO, P3CTI
, P3CTO, P3EI1, P3EI2, P3EI3, P3EI4, P3EI5, P3EI6, P3EI7, P3EI8, P3EL, P3ER, P3EO, P3RI, P3RL, P3RR, P3RO1, P3RO2, P3RO3, P3RO4, P3RO5, P3RO6
, P3RO7, P3RO8, P4CI1, P4CL, P4CR, P4CO, P4CTI, P4CTO, P4EI1, P4EI2, P4EI3, P4EI4, P4EI5, P4EI6, P4EI7, P4EI8, P4EL, P4ER, P4EO, P4RI, P4RL
, P4RR, P4RO1, P4RO2, P4RO3, P4RO4, P4RO5, P4RO6, P4RO7, P4RO8, P5CI1, P5CL, P5CR, P5CO, P5CTI, P5CTO, P5EI1, P5EI2, P5EI3, P5EI4, P5EI5, P5EI6
, P5EI7, P5EI8, P5EL, P5ER, P5EO, P5RI, P5RL, P5RR, P5RO1, P5RO2, P5RO3, P5RO4, P5RO5, P5RO6, P5RO7, P5RO8, P6CI1, P6CL, P6CR, P6CO, P6CTI
, P6CTO, P6EI1, P6EI2, P6EI3, P6EI4, P6EI5, P6EI6, P6EI7, P6EI8, P6EL, P6ER, P6EO, P6RI, P6RL, P6RR, P6RO1, P6RO2, P6RO3, P6RO4, P6RO5, P6RO6
, P6RO7, P6RO8, P7CI1, P7CL, P7CR, P7CO, P7CTI, P7CTO, P7EI1, P7EI2, P7EI3, P7EI4, P7EI5, P7EI6, P7EI7, P7EI8, P7EL, P7ER, P7EO, P7RI, P7RL
, P7RR, P7RO1, P7RO2, P7RO3, P7RO4, P7RO5, P7RO6, P7RO7, P7RO8, P8CI1, P8CL, P8CR, P8CO, P8CTI, P8CTO, P8EI1, P8EI2, P8EI3, P8EI4, P8EI5, P8EI6
, P8EI7, P8EI8, P8EL, P8ER, P8EO, P8RI, P8RL, P8RR, P8RO1, P8RO2, P8RO3, P8RO4, P8RO5, P8RO6, P8RO7, P8RO8, P9CI1, P9CL, P9CR, P9CO, P9CTI
, P9CTO, P9EI1, P9EI2, P9EI3, P9EI4, P9EI5, P9EI6, P9EI7, P9EI8, P9EL, P9ER, P9EO, P9RI, P9RL, P9RR, P9RO1, P9RO2, P9RO3, P9RO4, P9RO5, P9RO6
, P9RO7, P9RO8, P10CI1, P10CL, P10CR, P10CO, P10CTI, P10CTO, P10EI1, P10EI2, P10EI3, P10EI4, P10EI5, P10EI6, P10EI7, P10EI8, P10EL, P10ER, P10EO, P10RI, P10RL
, P10RR, P10RO1, P10RO2, P10RO3, P10RO4, P10RO5, P10RO6, P10RO7, P10RO8, P11CI1, P11CL, P11CR, P11CO, P11CTI, P11CTO, P11EI1, P11EI2, P11EI3, P11EI4, P11EI5, P11EI6
, P11EI7, P11EI8, P11EL, P11ER, P11EO, P11RI, P11RL, P11RR, P11RO1, P11RO2, P11RO3, P11RO4, P11RO5, P11RO6, P11RO7, P11RO8, P12CI1, P12CL, P12CR, P12CO, P12CTI
, P12CTO, P12EI1, P12EI2, P12EI3, P12EI4, P12EI5, P12EI6, P12EI7, P12EI8, P12EL, P12ER, P12EO, P12RI, P12RL, P12RR, P12RO1, P12RO2, P12RO3, P12RO4, P12RO5, P12RO6
, P12RO7, P12RO8, P13CI1, P13CL, P13CR, P13CO, P13CTI, P13CTO, P13EI1, P13EI2, P13EI3, P13EI4, P13EI5, P13EI6, P13EI7, P13EI8, P13EL, P13ER, P13EO, P13RI, P13RL
, P13RR, P13RO1, P13RO2, P13RO3, P13RO4, P13RO5, P13RO6, P13RO7, P13RO8, P14CI1, P14CL, P14CR, P14CO, P14CTI, P14CTO, P14EI1, P14EI2, P14EI3, P14EI4, P14EI5, P14EI6
, P14EI7, P14EI8, P14EL, P14ER, P14EO, P14RI, P14RL, P14RR, P14RO1, P14RO2, P14RO3, P14RO4, P14RO5, P14RO6, P14RO7, P14RO8, P15CI1, P15CL, P15CR, P15CO, P15CTI
, P15CTO, P15EI1, P15EI2, P15EI3, P15EI4, P15EI5, P15EI6, P15EI7, P15EI8, P15EL, P15ER, P15EO, P15RI, P15RL, P15RR, P15RO1, P15RO2, P15RO3, P15RO4, P15RO5, P15RO6
, P15RO7, P15RO8, P16CI1, P16CL, P16CR, P16CO, P16CTI, P16CTO, P16EI1, P16EI2, P16EI3, P16EI4, P16EI5, P16EI6, P16EI7, P16EI8, P16EL, P16ER, P16EO, P16RI, P16RL
, P16RR, P16RO1, P16RO2, P16RO3, P16RO4, P16RO5, P16RO6, P16RO7, P16RO8, P17CI1, P17CL, P17CR, P17CO, P17CTI, P17CTO, P17EI1, P17EI2, P17EI3, P17EI4, P17EI5, P17EI6
, P17EI7, P17EI8, P17EL, P17ER, P17EO, P17RI, P17RL, P17RR, P17RO1, P17RO2, P17RO3, P17RO4, P17RO5, P17RO6, P17RO7, P17RO8, P18CI1, P18CL, P18CR, P18CO, P18CTI
, P18CTO, P18EI1, P18EI2, P18EI3, P18EI4, P18EI5, P18EI6, P18EI7, P18EI8, P18EL, P18ER, P18EO, P18RI, P18RL, P18RR, P18RO1, P18RO2, P18RO3, P18RO4, P18RO5, P18RO6
, P18RO7, P18RO8, P19CI1, P19CL, P19CR, P19CO, P19CTI, P19CTO, P19EI1, P19EI2, P19EI3, P19EI4, P19EI5, P19EI6, P19EI7, P19EI8, P19EL, P19ER, P19EO, P19RI, P19RL
, P19RR, P19RO1, P19RO2, P19RO3, P19RO4, P19RO5, P19RO6, P19RO7, P19RO8, P20CI1, P20CL, P20CR, P20CO, P20CTI, P20CTO, P20EI1, P20EI2, P20EI3, P20EI4, P20EI5, P20EI6
, P20EI7, P20EI8, P20EL, P20ER, P20EO, P20RI, P20RL, P20RR, P20RO1, P20RO2, P20RO3, P20RO4, P20RO5, P20RO6, P20RO7, P20RO8, P21CI1, P21CL, P21CR, P21CO, P21CTI
, P21CTO, P21EI1, P21EI2, P21EI3, P21EI4, P21EI5, P21EI6, P21EI7, P21EI8, P21EL, P21ER, P21EO, P21RI, P21RL, P21RR, P21RO1, P21RO2, P21RO3, P21RO4, P21RO5, P21RO6
, P21RO7, P21RO8, P22CI1, P22CL, P22CR, P22CO, P22CTI, P22CTO, P22EI1, P22EI2, P22EI3, P22EI4, P22EI5, P22EI6, P22EI7, P22EI8, P22EL, P22ER, P22EO, P22RI, P22RL
, P22RR, P22RO1, P22RO2, P22RO3, P22RO4, P22RO5, P22RO6, P22RO7, P22RO8, P23CI1, P23CL, P23CR, P23CO, P23CTI, P23CTO, P23EI1, P23EI2, P23EI3, P23EI4, P23EI5, P23EI6
, P23EI7, P23EI8, P23EL, P23ER, P23EO, P23RI, P23RL, P23RR, P23RO1, P23RO2, P23RO3, P23RO4, P23RO5, P23RO6, P23RO7, P23RO8, P24CI1, P24CL, P24CR, P24CO, P24CTI
, P24CTO, P24EI1, P24EI2, P24EI3, P24EI4, P24EI5, P24EI6, P24EI7, P24EI8, P24EL, P24ER, P24EO, P24RI, P24RL, P24RR, P24RO1, P24RO2, P24RO3, P24RO4, P24RO5, P24RO6
, P24RO7, P24RO8, P25CI1, P25CL, P25CR, P25CO, P25CTI, P25CTO, P25EI1, P25EI2, P25EI3, P25EI4, P25EI5, P25EI6, P25EI7, P25EI8, P25EL, P25ER, P25EO, P25RI, P25RL
, P25RR, P25RO1, P25RO2, P25RO3, P25RO4, P25RO5, P25RO6, P25RO7, P25RO8, P26CI1, P26CL, P26CR, P26CO, P26CTI, P26CTO, P26EI1, P26EI2, P26EI3, P26EI4, P26EI5, P26EI6
, P26EI7, P26EI8, P26EL, P26ER, P26EO, P26RI, P26RL, P26RR, P26RO1, P26RO2, P26RO3, P26RO4, P26RO5, P26RO6, P26RO7, P26RO8, P27CI1, P27CL, P27CR, P27CO, P27CTI
, P27CTO, P27EI1, P27EI2, P27EI3, P27EI4, P27EI5, P27EI6, P27EI7, P27EI8, P27EL, P27ER, P27EO, P27RI, P27RL, P27RR, P27RO1, P27RO2, P27RO3, P27RO4, P27RO5, P27RO6
, P27RO7, P27RO8, P28CI1, P28CL, P28CR, P28CO, P28CTI, P28CTO, P28EI1, P28EI2, P28EI3, P28EI4, P28EI5, P28EI6, P28EI7, P28EI8, P28EL, P28ER, P28EO, P28RI, P28RL
, P28RR, P28RO1, P28RO2, P28RO3, P28RO4, P28RO5, P28RO6, P28RO7, P28RO8, P29CI1, P29CL, P29CR, P29CO, P29CTI, P29CTO, P29EI1, P29EI2, P29EI3, P29EI4, P29EI5, P29EI6
, P29EI7, P29EI8, P29EL, P29ER, P29EO, P29RI, P29RL, P29RR, P29RO1, P29RO2, P29RO3, P29RO4, P29RO5, P29RO6, P29RO7, P29RO8, P30CI1, P30CL, P30CR, P30CO, P30CTI
, P30CTO, P30EI1, P30EI2, P30EI3, P30EI4, P30EI5, P30EI6, P30EI7, P30EI8, P30EL, P30ER, P30EO, P30RI, P30RL, P30RR, P30RO1, P30RO2, P30RO3, P30RO4, P30RO5, P30RO6
, P30RO7, P30RO8, P31CI1, P31CL, P31CR, P31CO, P31CTI, P31CTO, P31EI1, P31EI2, P31EI3, P31EI4, P31EI5, P31EI6, P31EI7, P31EI8, P31EL, P31ER, P31EO, P31RI, P31RL
, P31RR, P31RO1, P31RO2, P31RO3, P31RO4, P31RO5, P31RO6, P31RO7, P31RO8, P32CI1, P32CL, P32CR, P32CO, P32CTI, P32CTO, P32EI1, P32EI2, P32EI3, P32EI4, P32EI5, P32EI6
, P32EI7, P32EI8, P32EL, P32ER, P32EO, P32RI, P32RL, P32RR, P32RO1, P32RO2, P32RO3, P32RO4, P32RO5, P32RO6, P32RO7, P32RO8, P33CI1, P33CL, P33CR, P33CO, P33CTI
, P33CTO, P33EI1, P33EI2, P33EI3, P33EI4, P33EI5, P33EI6, P33EI7, P33EI8, P33EL, P33ER, P33EO, P33RI, P33RL, P33RR, P33RO1, P33RO2, P33RO3, P33RO4, P33RO5, P33RO6
, P33RO7, P33RO8, P34CI1, P34CL, P34CR, P34CO, P34CTI, P34CTO, P34EI1, P34EI2, P34EI3, P34EI4, P34EI5, P34EI6, P34EI7, P34EI8, P34EL, P34ER, P34EO, P34RI, P34RL
, P34RR, P34RO1, P34RO2, P34RO3, P34RO4, P34RO5, P34RO6, P34RO7, P34RO8);
    output AL1D;
    output AL1T;
    output AL2D;
    output AL2T;
    output AL3D;
    output AL3T;
    input ALCK1;
    input ALCK2;
    input ALCK3;
    input CA1D1;
    input CA1D2;
    input CA1D3;
    input CA1D4;
    input CA1D5;
    input CA1D6;
    input CA1N1;
    input CA1N2;
    input CA1N3;
    input CA1N4;
    input CA1P1;
    input CA1P2;
    input CA1P3;
    input CA1P4;
    input CA1T1;
    input CA1T2;
    input CA1T3;
    input CA1T4;
    input CA2D1;
    input CA2D2;
    input CA2D3;
    input CA2D4;
    input CA2D5;
    input CA2D6;
    input CA2N1;
    input CA2N2;
    input CA2N3;
    input CA2N4;
    input CA2P1;
    input CA2P2;
    input CA2P3;
    input CA2P4;
    input CA2T1;
    input CA2T2;
    input CA2T3;
    input CA2T4;
    input CCK;
    output CKO1;
    output CKO2;
    output DCL;
    input DCRN;
    input DQ1CI1;
    input DQ1CI2;
    input DQ1CI3;
    input DQ1CI4;
    input DQ1CI5;
    input DQ1CI6;
    input DQ1CI7;
    input DQ1CI8;
    input DQ2CI1;
    input DQ2CI2;
    input DQ2CI3;
    input DQ2CI4;
    input DQ2CI5;
    input DQ2CI6;
    input DQ2CI7;
    input DQ2CI8;
    input DQ3CI1;
    input DQ3CI2;
    input DQ3CI3;
    input DQ3CI4;
    input DQ3CI5;
    input DQ3CI6;
    input DQ3CI7;
    input DQ3CI8;
    input DQS1CI1;
    input DQS1CI2;
    input DQS1CI3;
    input DQS1CI4;
    input DQS1CI5;
    input DQS1CI6;
    input DQS1CI7;
    input DQS1CI8;
    input DQS2CI1;
    input DQS2CI2;
    input DQS2CI3;
    input DQS2CI4;
    input DQS2CI5;
    input DQS2CI6;
    input DQS2CI7;
    input DQS2CI8;
    input DQS3CI1;
    input DQS3CI2;
    input DQS3CI3;
    input DQS3CI4;
    input DQS3CI5;
    input DQS3CI6;
    input DQS3CI7;
    input DQS3CI8;
    input DRA1;
    input DRA2;
    input DRA3;
    input DRA4;
    input DRCCSN;
    input DRDPA1CSN;
    input DRDPA2CSN;
    input DRDPA3CSN;
    input DRE;
    input DRI1;
    input DRI1CSN;
    input DRI2;
    input DRI2CSN;
    input DRI3;
    input DRI3CSN;
    input DRI4;
    input DRI5;
    input DRI6;
    output DRO1;
    input DRO1CSN;
    output DRO2;
    input DRO2CSN;
    output DRO3;
    input DRO3CSN;
    output DRO4;
    output DRO5;
    output DRO6;
    input DRWDS;
    input DRWEN;
    input FA1;
    input FA2;
    input FA3;
    input FA4;
    input FA5;
    input FA6;
    input FCK1;
    input FCK2;
    input FDCK;
    output FLD;
    output FLG;
    input FZ;
    input LD1RN;
    input LD2RN;
    input LD3RN;
    input LDSCK1;
    input LDSCK2;
    input LDSCK3;
    input LE;
    input P10CI1;
    input P10CL;
    output P10CO;
    input P10CR;
    input P10CTI;
    output P10CTO;
    input P10EI1;
    input P10EI2;
    input P10EI3;
    input P10EI4;
    input P10EI5;
    input P10EI6;
    input P10EI7;
    input P10EI8;
    input P10EL;
    output P10EO;
    input P10ER;
    input P10RI;
    input P10RL;
    output P10RO1;
    output P10RO2;
    output P10RO3;
    output P10RO4;
    output P10RO5;
    output P10RO6;
    output P10RO7;
    output P10RO8;
    input P10RR;
    input P11CI1;
    input P11CL;
    output P11CO;
    input P11CR;
    input P11CTI;
    output P11CTO;
    input P11EI1;
    input P11EI2;
    input P11EI3;
    input P11EI4;
    input P11EI5;
    input P11EI6;
    input P11EI7;
    input P11EI8;
    input P11EL;
    output P11EO;
    input P11ER;
    input P11RI;
    input P11RL;
    output P11RO1;
    output P11RO2;
    output P11RO3;
    output P11RO4;
    output P11RO5;
    output P11RO6;
    output P11RO7;
    output P11RO8;
    input P11RR;
    input P12CI1;
    input P12CL;
    output P12CO;
    input P12CR;
    input P12CTI;
    output P12CTO;
    input P12EI1;
    input P12EI2;
    input P12EI3;
    input P12EI4;
    input P12EI5;
    input P12EI6;
    input P12EI7;
    input P12EI8;
    input P12EL;
    output P12EO;
    input P12ER;
    input P12RI;
    input P12RL;
    output P12RO1;
    output P12RO2;
    output P12RO3;
    output P12RO4;
    output P12RO5;
    output P12RO6;
    output P12RO7;
    output P12RO8;
    input P12RR;
    input P13CI1;
    input P13CL;
    output P13CO;
    input P13CR;
    input P13CTI;
    output P13CTO;
    input P13EI1;
    input P13EI2;
    input P13EI3;
    input P13EI4;
    input P13EI5;
    input P13EI6;
    input P13EI7;
    input P13EI8;
    input P13EL;
    output P13EO;
    input P13ER;
    input P13RI;
    input P13RL;
    output P13RO1;
    output P13RO2;
    output P13RO3;
    output P13RO4;
    output P13RO5;
    output P13RO6;
    output P13RO7;
    output P13RO8;
    input P13RR;
    input P14CI1;
    input P14CL;
    output P14CO;
    input P14CR;
    input P14CTI;
    output P14CTO;
    input P14EI1;
    input P14EI2;
    input P14EI3;
    input P14EI4;
    input P14EI5;
    input P14EI6;
    input P14EI7;
    input P14EI8;
    input P14EL;
    output P14EO;
    input P14ER;
    input P14RI;
    input P14RL;
    output P14RO1;
    output P14RO2;
    output P14RO3;
    output P14RO4;
    output P14RO5;
    output P14RO6;
    output P14RO7;
    output P14RO8;
    input P14RR;
    input P15CI1;
    input P15CL;
    output P15CO;
    input P15CR;
    input P15CTI;
    output P15CTO;
    input P15EI1;
    input P15EI2;
    input P15EI3;
    input P15EI4;
    input P15EI5;
    input P15EI6;
    input P15EI7;
    input P15EI8;
    input P15EL;
    output P15EO;
    input P15ER;
    input P15RI;
    input P15RL;
    output P15RO1;
    output P15RO2;
    output P15RO3;
    output P15RO4;
    output P15RO5;
    output P15RO6;
    output P15RO7;
    output P15RO8;
    input P15RR;
    input P16CI1;
    input P16CL;
    output P16CO;
    input P16CR;
    input P16CTI;
    output P16CTO;
    input P16EI1;
    input P16EI2;
    input P16EI3;
    input P16EI4;
    input P16EI5;
    input P16EI6;
    input P16EI7;
    input P16EI8;
    input P16EL;
    output P16EO;
    input P16ER;
    input P16RI;
    input P16RL;
    output P16RO1;
    output P16RO2;
    output P16RO3;
    output P16RO4;
    output P16RO5;
    output P16RO6;
    output P16RO7;
    output P16RO8;
    input P16RR;
    input P17CI1;
    input P17CL;
    output P17CO;
    input P17CR;
    input P17CTI;
    output P17CTO;
    input P17EI1;
    input P17EI2;
    input P17EI3;
    input P17EI4;
    input P17EI5;
    input P17EI6;
    input P17EI7;
    input P17EI8;
    input P17EL;
    output P17EO;
    input P17ER;
    input P17RI;
    input P17RL;
    output P17RO1;
    output P17RO2;
    output P17RO3;
    output P17RO4;
    output P17RO5;
    output P17RO6;
    output P17RO7;
    output P17RO8;
    input P17RR;
    input P18CI1;
    input P18CL;
    output P18CO;
    input P18CR;
    input P18CTI;
    output P18CTO;
    input P18EI1;
    input P18EI2;
    input P18EI3;
    input P18EI4;
    input P18EI5;
    input P18EI6;
    input P18EI7;
    input P18EI8;
    input P18EL;
    output P18EO;
    input P18ER;
    input P18RI;
    input P18RL;
    output P18RO1;
    output P18RO2;
    output P18RO3;
    output P18RO4;
    output P18RO5;
    output P18RO6;
    output P18RO7;
    output P18RO8;
    input P18RR;
    input P19CI1;
    input P19CL;
    output P19CO;
    input P19CR;
    input P19CTI;
    output P19CTO;
    input P19EI1;
    input P19EI2;
    input P19EI3;
    input P19EI4;
    input P19EI5;
    input P19EI6;
    input P19EI7;
    input P19EI8;
    input P19EL;
    output P19EO;
    input P19ER;
    input P19RI;
    input P19RL;
    output P19RO1;
    output P19RO2;
    output P19RO3;
    output P19RO4;
    output P19RO5;
    output P19RO6;
    output P19RO7;
    output P19RO8;
    input P19RR;
    input P1CI1;
    input P1CL;
    output P1CO;
    input P1CR;
    input P1CTI;
    output P1CTO;
    input P1EI1;
    input P1EI2;
    input P1EI3;
    input P1EI4;
    input P1EI5;
    input P1EI6;
    input P1EI7;
    input P1EI8;
    input P1EL;
    output P1EO;
    input P1ER;
    input P1RI;
    input P1RL;
    output P1RO1;
    output P1RO2;
    output P1RO3;
    output P1RO4;
    output P1RO5;
    output P1RO6;
    output P1RO7;
    output P1RO8;
    input P1RR;
    input P20CI1;
    input P20CL;
    output P20CO;
    input P20CR;
    input P20CTI;
    output P20CTO;
    input P20EI1;
    input P20EI2;
    input P20EI3;
    input P20EI4;
    input P20EI5;
    input P20EI6;
    input P20EI7;
    input P20EI8;
    input P20EL;
    output P20EO;
    input P20ER;
    input P20RI;
    input P20RL;
    output P20RO1;
    output P20RO2;
    output P20RO3;
    output P20RO4;
    output P20RO5;
    output P20RO6;
    output P20RO7;
    output P20RO8;
    input P20RR;
    input P21CI1;
    input P21CL;
    output P21CO;
    input P21CR;
    input P21CTI;
    output P21CTO;
    input P21EI1;
    input P21EI2;
    input P21EI3;
    input P21EI4;
    input P21EI5;
    input P21EI6;
    input P21EI7;
    input P21EI8;
    input P21EL;
    output P21EO;
    input P21ER;
    input P21RI;
    input P21RL;
    output P21RO1;
    output P21RO2;
    output P21RO3;
    output P21RO4;
    output P21RO5;
    output P21RO6;
    output P21RO7;
    output P21RO8;
    input P21RR;
    input P22CI1;
    input P22CL;
    output P22CO;
    input P22CR;
    input P22CTI;
    output P22CTO;
    input P22EI1;
    input P22EI2;
    input P22EI3;
    input P22EI4;
    input P22EI5;
    input P22EI6;
    input P22EI7;
    input P22EI8;
    input P22EL;
    output P22EO;
    input P22ER;
    input P22RI;
    input P22RL;
    output P22RO1;
    output P22RO2;
    output P22RO3;
    output P22RO4;
    output P22RO5;
    output P22RO6;
    output P22RO7;
    output P22RO8;
    input P22RR;
    input P23CI1;
    input P23CL;
    output P23CO;
    input P23CR;
    input P23CTI;
    output P23CTO;
    input P23EI1;
    input P23EI2;
    input P23EI3;
    input P23EI4;
    input P23EI5;
    input P23EI6;
    input P23EI7;
    input P23EI8;
    input P23EL;
    output P23EO;
    input P23ER;
    input P23RI;
    input P23RL;
    output P23RO1;
    output P23RO2;
    output P23RO3;
    output P23RO4;
    output P23RO5;
    output P23RO6;
    output P23RO7;
    output P23RO8;
    input P23RR;
    input P24CI1;
    input P24CL;
    output P24CO;
    input P24CR;
    input P24CTI;
    output P24CTO;
    input P24EI1;
    input P24EI2;
    input P24EI3;
    input P24EI4;
    input P24EI5;
    input P24EI6;
    input P24EI7;
    input P24EI8;
    input P24EL;
    output P24EO;
    input P24ER;
    input P24RI;
    input P24RL;
    output P24RO1;
    output P24RO2;
    output P24RO3;
    output P24RO4;
    output P24RO5;
    output P24RO6;
    output P24RO7;
    output P24RO8;
    input P24RR;
    input P25CI1;
    input P25CL;
    output P25CO;
    input P25CR;
    input P25CTI;
    output P25CTO;
    input P25EI1;
    input P25EI2;
    input P25EI3;
    input P25EI4;
    input P25EI5;
    input P25EI6;
    input P25EI7;
    input P25EI8;
    input P25EL;
    output P25EO;
    input P25ER;
    input P25RI;
    input P25RL;
    output P25RO1;
    output P25RO2;
    output P25RO3;
    output P25RO4;
    output P25RO5;
    output P25RO6;
    output P25RO7;
    output P25RO8;
    input P25RR;
    input P26CI1;
    input P26CL;
    output P26CO;
    input P26CR;
    input P26CTI;
    output P26CTO;
    input P26EI1;
    input P26EI2;
    input P26EI3;
    input P26EI4;
    input P26EI5;
    input P26EI6;
    input P26EI7;
    input P26EI8;
    input P26EL;
    output P26EO;
    input P26ER;
    input P26RI;
    input P26RL;
    output P26RO1;
    output P26RO2;
    output P26RO3;
    output P26RO4;
    output P26RO5;
    output P26RO6;
    output P26RO7;
    output P26RO8;
    input P26RR;
    input P27CI1;
    input P27CL;
    output P27CO;
    input P27CR;
    input P27CTI;
    output P27CTO;
    input P27EI1;
    input P27EI2;
    input P27EI3;
    input P27EI4;
    input P27EI5;
    input P27EI6;
    input P27EI7;
    input P27EI8;
    input P27EL;
    output P27EO;
    input P27ER;
    input P27RI;
    input P27RL;
    output P27RO1;
    output P27RO2;
    output P27RO3;
    output P27RO4;
    output P27RO5;
    output P27RO6;
    output P27RO7;
    output P27RO8;
    input P27RR;
    input P28CI1;
    input P28CL;
    output P28CO;
    input P28CR;
    input P28CTI;
    output P28CTO;
    input P28EI1;
    input P28EI2;
    input P28EI3;
    input P28EI4;
    input P28EI5;
    input P28EI6;
    input P28EI7;
    input P28EI8;
    input P28EL;
    output P28EO;
    input P28ER;
    input P28RI;
    input P28RL;
    output P28RO1;
    output P28RO2;
    output P28RO3;
    output P28RO4;
    output P28RO5;
    output P28RO6;
    output P28RO7;
    output P28RO8;
    input P28RR;
    input P29CI1;
    input P29CL;
    output P29CO;
    input P29CR;
    input P29CTI;
    output P29CTO;
    input P29EI1;
    input P29EI2;
    input P29EI3;
    input P29EI4;
    input P29EI5;
    input P29EI6;
    input P29EI7;
    input P29EI8;
    input P29EL;
    output P29EO;
    input P29ER;
    input P29RI;
    input P29RL;
    output P29RO1;
    output P29RO2;
    output P29RO3;
    output P29RO4;
    output P29RO5;
    output P29RO6;
    output P29RO7;
    output P29RO8;
    input P29RR;
    input P2CI1;
    input P2CL;
    output P2CO;
    input P2CR;
    input P2CTI;
    output P2CTO;
    input P2EI1;
    input P2EI2;
    input P2EI3;
    input P2EI4;
    input P2EI5;
    input P2EI6;
    input P2EI7;
    input P2EI8;
    input P2EL;
    output P2EO;
    input P2ER;
    input P2RI;
    input P2RL;
    output P2RO1;
    output P2RO2;
    output P2RO3;
    output P2RO4;
    output P2RO5;
    output P2RO6;
    output P2RO7;
    output P2RO8;
    input P2RR;
    input P30CI1;
    input P30CL;
    output P30CO;
    input P30CR;
    input P30CTI;
    output P30CTO;
    input P30EI1;
    input P30EI2;
    input P30EI3;
    input P30EI4;
    input P30EI5;
    input P30EI6;
    input P30EI7;
    input P30EI8;
    input P30EL;
    output P30EO;
    input P30ER;
    input P30RI;
    input P30RL;
    output P30RO1;
    output P30RO2;
    output P30RO3;
    output P30RO4;
    output P30RO5;
    output P30RO6;
    output P30RO7;
    output P30RO8;
    input P30RR;
    input P31CI1;
    input P31CL;
    output P31CO;
    input P31CR;
    input P31CTI;
    output P31CTO;
    input P31EI1;
    input P31EI2;
    input P31EI3;
    input P31EI4;
    input P31EI5;
    input P31EI6;
    input P31EI7;
    input P31EI8;
    input P31EL;
    output P31EO;
    input P31ER;
    input P31RI;
    input P31RL;
    output P31RO1;
    output P31RO2;
    output P31RO3;
    output P31RO4;
    output P31RO5;
    output P31RO6;
    output P31RO7;
    output P31RO8;
    input P31RR;
    input P32CI1;
    input P32CL;
    output P32CO;
    input P32CR;
    input P32CTI;
    output P32CTO;
    input P32EI1;
    input P32EI2;
    input P32EI3;
    input P32EI4;
    input P32EI5;
    input P32EI6;
    input P32EI7;
    input P32EI8;
    input P32EL;
    output P32EO;
    input P32ER;
    input P32RI;
    input P32RL;
    output P32RO1;
    output P32RO2;
    output P32RO3;
    output P32RO4;
    output P32RO5;
    output P32RO6;
    output P32RO7;
    output P32RO8;
    input P32RR;
    input P33CI1;
    input P33CL;
    output P33CO;
    input P33CR;
    input P33CTI;
    output P33CTO;
    input P33EI1;
    input P33EI2;
    input P33EI3;
    input P33EI4;
    input P33EI5;
    input P33EI6;
    input P33EI7;
    input P33EI8;
    input P33EL;
    output P33EO;
    input P33ER;
    input P33RI;
    input P33RL;
    output P33RO1;
    output P33RO2;
    output P33RO3;
    output P33RO4;
    output P33RO5;
    output P33RO6;
    output P33RO7;
    output P33RO8;
    input P33RR;
    input P34CI1;
    input P34CL;
    output P34CO;
    input P34CR;
    input P34CTI;
    output P34CTO;
    input P34EI1;
    input P34EI2;
    input P34EI3;
    input P34EI4;
    input P34EI5;
    input P34EI6;
    input P34EI7;
    input P34EI8;
    input P34EL;
    output P34EO;
    input P34ER;
    input P34RI;
    input P34RL;
    output P34RO1;
    output P34RO2;
    output P34RO3;
    output P34RO4;
    output P34RO5;
    output P34RO6;
    output P34RO7;
    output P34RO8;
    input P34RR;
    input P3CI1;
    input P3CL;
    output P3CO;
    input P3CR;
    input P3CTI;
    output P3CTO;
    input P3EI1;
    input P3EI2;
    input P3EI3;
    input P3EI4;
    input P3EI5;
    input P3EI6;
    input P3EI7;
    input P3EI8;
    input P3EL;
    output P3EO;
    input P3ER;
    input P3RI;
    input P3RL;
    output P3RO1;
    output P3RO2;
    output P3RO3;
    output P3RO4;
    output P3RO5;
    output P3RO6;
    output P3RO7;
    output P3RO8;
    input P3RR;
    input P4CI1;
    input P4CL;
    output P4CO;
    input P4CR;
    input P4CTI;
    output P4CTO;
    input P4EI1;
    input P4EI2;
    input P4EI3;
    input P4EI4;
    input P4EI5;
    input P4EI6;
    input P4EI7;
    input P4EI8;
    input P4EL;
    output P4EO;
    input P4ER;
    input P4RI;
    input P4RL;
    output P4RO1;
    output P4RO2;
    output P4RO3;
    output P4RO4;
    output P4RO5;
    output P4RO6;
    output P4RO7;
    output P4RO8;
    input P4RR;
    input P5CI1;
    input P5CL;
    output P5CO;
    input P5CR;
    input P5CTI;
    output P5CTO;
    input P5EI1;
    input P5EI2;
    input P5EI3;
    input P5EI4;
    input P5EI5;
    input P5EI6;
    input P5EI7;
    input P5EI8;
    input P5EL;
    output P5EO;
    input P5ER;
    input P5RI;
    input P5RL;
    output P5RO1;
    output P5RO2;
    output P5RO3;
    output P5RO4;
    output P5RO5;
    output P5RO6;
    output P5RO7;
    output P5RO8;
    input P5RR;
    input P6CI1;
    input P6CL;
    output P6CO;
    input P6CR;
    input P6CTI;
    output P6CTO;
    input P6EI1;
    input P6EI2;
    input P6EI3;
    input P6EI4;
    input P6EI5;
    input P6EI6;
    input P6EI7;
    input P6EI8;
    input P6EL;
    output P6EO;
    input P6ER;
    input P6RI;
    input P6RL;
    output P6RO1;
    output P6RO2;
    output P6RO3;
    output P6RO4;
    output P6RO5;
    output P6RO6;
    output P6RO7;
    output P6RO8;
    input P6RR;
    input P7CI1;
    input P7CL;
    output P7CO;
    input P7CR;
    input P7CTI;
    output P7CTO;
    input P7EI1;
    input P7EI2;
    input P7EI3;
    input P7EI4;
    input P7EI5;
    input P7EI6;
    input P7EI7;
    input P7EI8;
    input P7EL;
    output P7EO;
    input P7ER;
    input P7RI;
    input P7RL;
    output P7RO1;
    output P7RO2;
    output P7RO3;
    output P7RO4;
    output P7RO5;
    output P7RO6;
    output P7RO7;
    output P7RO8;
    input P7RR;
    input P8CI1;
    input P8CL;
    output P8CO;
    input P8CR;
    input P8CTI;
    output P8CTO;
    input P8EI1;
    input P8EI2;
    input P8EI3;
    input P8EI4;
    input P8EI5;
    input P8EI6;
    input P8EI7;
    input P8EI8;
    input P8EL;
    output P8EO;
    input P8ER;
    input P8RI;
    input P8RL;
    output P8RO1;
    output P8RO2;
    output P8RO3;
    output P8RO4;
    output P8RO5;
    output P8RO6;
    output P8RO7;
    output P8RO8;
    input P8RR;
    input P9CI1;
    input P9CL;
    output P9CO;
    input P9CR;
    input P9CTI;
    output P9CTO;
    input P9EI1;
    input P9EI2;
    input P9EI3;
    input P9EI4;
    input P9EI5;
    input P9EI6;
    input P9EI7;
    input P9EI8;
    input P9EL;
    output P9EO;
    input P9ER;
    input P9RI;
    input P9RL;
    output P9RO1;
    output P9RO2;
    output P9RO3;
    output P9RO4;
    output P9RO5;
    output P9RO6;
    output P9RO7;
    output P9RO8;
    input P9RR;
    input SE;
    input SWRX1CK;
    input SWRX2CK;
    parameter cal_delay1 = "";
    parameter cal_delay2 = "";
    parameter div1 = 3'b000;
    parameter div2 = 3'b000;
    parameter div3 = 3'b000;
    parameter div_swrx1 = 3'b000;
    parameter div_swrx2 = 3'b000;
    parameter inv_ld_sck1 = 1'b0;
    parameter inv_ld_sck2 = 1'b0;
    parameter inv_ld_sck3 = 1'b0;
    parameter link_ld_12 = 1'b0;
    parameter link_ld_23 = 1'b0;
    parameter mode_side1 = 0;
    parameter mode_side2 = 0;
    parameter mode_side3 = 0;
    parameter pads_dict = "";
    parameter pads_path = "";
    parameter sel_clk_out1 = 1'b0;
    parameter sel_clk_out2 = 1'b0;
    parameter sel_dc_clk = 2'b00;
    parameter sel_ld_fck1 = 2'b00;
    parameter sel_ld_fck2 = 2'b00;
    parameter sel_ld_fck3 = 2'b00;
    parameter sel_sw_fck1 = 2'b00;
    parameter sel_sw_fck2 = 2'b00;
    parameter use_dc = 1'b0;
endmodule

//(* blackbox *)
//module NX_LUT(I1, I2, I3, I4, O);
//    input I1;
//    input I2;
//    input I3;
//    input I4;
//    output O;
//    parameter lut_table = 16'b0000000000000000;
//endmodule

(* blackbox *)
module NX_PLL(REF, FBK, VCO, D1, D2, D3, OSC, RDY);
    output D1;
    output D2;
    output D3;
    input FBK;
    output OSC;
    output RDY;
    input REF;
    output VCO;
    parameter clk_outdiv1 = 0;
    parameter clk_outdiv2 = 0;
    parameter clk_outdiv3 = 0;
    parameter ext_fbk_on = 1'b0;
    parameter fbk_delay = 0;
    parameter fbk_delay_on = 1'b0;
    parameter fbk_div_on = 1'b0;
    parameter fbk_intdiv = 2;
    parameter location = "";
    parameter ref_div_on = 1'b0;
    parameter vco_range = 0;
endmodule

(* blackbox *)
module NX_PLL_L(REF, FBK, R, VCO, LDFO, REFO, DIVO1, DIVO2, DIVP1, DIVP2, DIVP3, OSC, PLL_LOCKED, CAL_LOCKED);
    output CAL_LOCKED;
    output DIVO1;
    output DIVO2;
    output DIVP1;
    output DIVP2;
    output DIVP3;
    input FBK;
    output LDFO;
    output OSC;
    output PLL_LOCKED;
    input R;
    input REF;
    output REFO;
    output VCO;
    parameter cfg_use_pll = 1'b1;
    parameter clk_outdivo1 = 0;
    parameter clk_outdivp1 = 0;
    parameter clk_outdivp2 = 0;
    parameter clk_outdivp3o2 = 0;
    parameter ext_fbk_on = 1'b0;
    parameter fbk_delay = 0;
    parameter fbk_delay_on = 1'b0;
    parameter fbk_intdiv = 2;
    parameter location = "";
    parameter pll_cpump = 3'b010;
    parameter ref_intdiv = 0;
    parameter ref_osc_on = 1'b0;
    parameter wfg_sync_cal_lock = 1'b0;
    parameter wfg_sync_pll_lock = 1'b0;
endmodule

(* blackbox *)
module NX_PLL_U(R, REF, FBK, OSC, VCO, LDFO, REFO, CLK_DIV1, CLK_DIV2, CLK_DIV3, CLK_DIV4, CLK_DIVD1, CLK_DIVD2, CLK_DIVD3, CLK_DIVD4, CLK_DIVD5, PLL_LOCKED, PLL_LOCKEDA, ARST_CAL, CLK_CAL, CLK_CAL_DIV
, CAL_LOCKED, EXT_CAL_LOCKED, CAL1, CAL2, CAL3, CAL4, CAL5, EXT_CAL1, EXT_CAL2, EXT_CAL3, EXT_CAL4, EXT_CAL5);
    input ARST_CAL;
    output CAL1;
    output CAL2;
    output CAL3;
    output CAL4;
    output CAL5;
    output CAL_LOCKED;
    input CLK_CAL;
    output CLK_CAL_DIV;
    output CLK_DIV1;
    output CLK_DIV2;
    output CLK_DIV3;
    output CLK_DIV4;
    output CLK_DIVD1;
    output CLK_DIVD2;
    output CLK_DIVD3;
    output CLK_DIVD4;
    output CLK_DIVD5;
    input EXT_CAL1;
    input EXT_CAL2;
    input EXT_CAL3;
    input EXT_CAL4;
    input EXT_CAL5;
    input EXT_CAL_LOCKED;
    input FBK;
    output LDFO;
    output OSC;
    output PLL_LOCKED;
    output PLL_LOCKEDA;
    input R;
    input REF;
    output REFO;
    output VCO;
    parameter cal_delay = 6'b011011;
    parameter cal_div = 4'b0111;
    parameter clk_cal_sel = 2'b01;
    parameter clk_outdiv1 = 3'b000;
    parameter clk_outdiv2 = 3'b000;
    parameter clk_outdiv3 = 3'b000;
    parameter clk_outdiv4 = 3'b000;
    parameter clk_outdivd1 = 4'b0000;
    parameter clk_outdivd2 = 4'b0000;
    parameter clk_outdivd3 = 4'b0000;
    parameter clk_outdivd4 = 4'b0000;
    parameter clk_outdivd5 = 4'b0000;
    parameter ext_fbk_on = 1'b0;
    parameter fbk_delay = 6'b000000;
    parameter fbk_delay_on = 1'b0;
    parameter fbk_intdiv = 7'b0000000;
    parameter location = "";
    parameter pll_cpump = 4'b0000;
    parameter pll_lock = 4'b0000;
    parameter pll_lpf_cap = 4'b0000;
    parameter pll_lpf_res = 4'b0000;
    parameter pll_odf = 2'b00;
    parameter ref_intdiv = 5'b00000;
    parameter ref_osc_on = 1'b0;
    parameter use_cal = 1'b0;
    parameter use_pll = 1'b1;
endmodule

(* blackbox *)
module NX_PLL_U_WRAP(R, REF, FBK, OSC, VCO, LDFO, REFO, PLL_LOCKED, PLL_LOCKEDA, ARST_CAL, CLK_CAL, CLK_CAL_DIV, CAL_LOCKED, EXT_CAL_LOCKED, CAL, CLK_DIVD, EXT_CAL, CLK_DIV);
    input ARST_CAL;
    output [4:0] CAL;
    output CAL_LOCKED;
    input CLK_CAL;
    output CLK_CAL_DIV;
    output [3:0] CLK_DIV;
    output [4:0] CLK_DIVD;
    input [4:0] EXT_CAL;
    input EXT_CAL_LOCKED;
    input FBK;
    output LDFO;
    output OSC;
    output PLL_LOCKED;
    output PLL_LOCKEDA;
    input R;
    input REF;
    output REFO;
    output VCO;
    parameter cal_delay = 6'b011011;
    parameter cal_div = 4'b0111;
    parameter clk_cal_sel = 2'b01;
    parameter clk_outdiv1 = 3'b000;
    parameter clk_outdiv2 = 3'b000;
    parameter clk_outdiv3 = 3'b000;
    parameter clk_outdiv4 = 3'b000;
    parameter clk_outdivd1 = 4'b0000;
    parameter clk_outdivd2 = 4'b0000;
    parameter clk_outdivd3 = 4'b0000;
    parameter clk_outdivd4 = 4'b0000;
    parameter clk_outdivd5 = 4'b0000;
    parameter ext_fbk_on = 1'b0;
    parameter fbk_delay = 6'b000000;
    parameter fbk_delay_on = 1'b0;
    parameter fbk_intdiv = 7'b0000000;
    parameter location = "";
    parameter pll_cpump = 4'b0000;
    parameter pll_lock = 4'b0000;
    parameter pll_lpf_cap = 4'b0000;
    parameter pll_lpf_res = 4'b0000;
    parameter pll_odf = 2'b00;
    parameter ref_intdiv = 5'b00000;
    parameter ref_osc_on = 1'b0;
    parameter use_cal = 1'b0;
    parameter use_pll = 1'b1;
endmodule

(* blackbox *)
module NX_PMA_L(CLK_USER_I, CLK_REF_I, PRE_SG_I, PRE_EN_I, PRE_IS_I1, PRE_IS_I2, PRE_IS_I3, PRE_IS_I4, MAIN_SG_I, MAIN_EN_I1, MAIN_EN_I2, MAIN_EN_I3, MAIN_EN_I4, MAIN_EN_I5, MAIN_EN_I6, MARG_S_I1, MARG_S_I2, MARG_S_I3, MARG_S_I4, MARG_IS_I1, MARG_IS_I2
, MARG_IS_I3, MARG_IS_I4, MARG_SV_I1, MARG_SV_I2, MARG_SV_I3, MARG_SV_I4, MARG_SV_I5, MARG_ISV_I1, MARG_ISV_I2, MARG_ISV_I3, MARG_ISV_I4, MARG_ISV_I5, POST_EN_I1, POST_EN_I2, POST_EN_I3, POST_EN_I4, POST_EN_I5, POST_SG_I, POST_IS_I1, POST_IS_I2, POST_IS_I3
, POST_IS_I4, POST_ISV_I1, POST_ISV_I2, POST_ISV_I3, POST_ISV_I4, TX_SEL_I1, TX_SEL_I2, TX_SEL_I3, TX_SEL_I4, TX_SEL_I5, TX_SEL_I6, CT_CAP_I1, CT_CAP_I2, CT_CAP_I3, CT_CAP_I4, CT_RESP_I1, CT_RESP_I2, CT_RESP_I3, CT_RESP_I4, CT_RESN_I1, CT_RESN_I2
, CT_RESN_I3, CT_RESN_I4, M_EYE_I, RX_SEL_I1, RX_SEL_I2, RX_SEL_I3, RX_SEL_I4, RX_SEL_I5, RX_SEL_I6, PLL_RN_I, RST_N_I, CAL_1P_I1, CAL_1P_I2, CAL_1P_I3, CAL_1P_I4, CAL_1P_I5, CAL_1P_I6, CAL_1P_I7, CAL_1P_I8, CAL_2N_I1, CAL_2N_I2
, CAL_2N_I3, CAL_2N_I4, CAL_2N_I5, CAL_2N_I6, CAL_2N_I7, CAL_2N_I8, CAL_3N_I1, CAL_3N_I2, CAL_3N_I3, CAL_3N_I4, CAL_3N_I5, CAL_3N_I6, CAL_3N_I7, CAL_3N_I8, CAL_4P_I1, CAL_4P_I2, CAL_4P_I3, CAL_4P_I4, CAL_4P_I5, CAL_4P_I6, CAL_4P_I7
, CAL_4P_I8, CAL_SEL_I1, CAL_SEL_I2, CAL_SEL_I3, CAL_SEL_I4, CAL_E_I, LOCK_E_I, OVS_E_I, TST_I1, TST_I2, TST_I3, TST_I4, TST_I5, TST_I6, TST_I7, TST_I8, CLK_O, LOCK_O, CAL_O, TST_O1, TST_O2
, TST_O3, TST_O4, TST_O5, TST_O6, TST_O7, TST_O8, CLK_EXT_I, LINK_TX1, LINK_TX2, LINK_TX3, LINK_TX4, LINK_TX5, LINK_RX0, LINK_RX1, LINK_RX2, LINK_RX3, LINK_RX4, LINK_RX5, LINK_TX0);
    input CAL_1P_I1;
    input CAL_1P_I2;
    input CAL_1P_I3;
    input CAL_1P_I4;
    input CAL_1P_I5;
    input CAL_1P_I6;
    input CAL_1P_I7;
    input CAL_1P_I8;
    input CAL_2N_I1;
    input CAL_2N_I2;
    input CAL_2N_I3;
    input CAL_2N_I4;
    input CAL_2N_I5;
    input CAL_2N_I6;
    input CAL_2N_I7;
    input CAL_2N_I8;
    input CAL_3N_I1;
    input CAL_3N_I2;
    input CAL_3N_I3;
    input CAL_3N_I4;
    input CAL_3N_I5;
    input CAL_3N_I6;
    input CAL_3N_I7;
    input CAL_3N_I8;
    input CAL_4P_I1;
    input CAL_4P_I2;
    input CAL_4P_I3;
    input CAL_4P_I4;
    input CAL_4P_I5;
    input CAL_4P_I6;
    input CAL_4P_I7;
    input CAL_4P_I8;
    input CAL_E_I;
    output CAL_O;
    input CAL_SEL_I1;
    input CAL_SEL_I2;
    input CAL_SEL_I3;
    input CAL_SEL_I4;
    input CLK_EXT_I;
    output CLK_O;
    input CLK_REF_I;
    input CLK_USER_I;
    input CT_CAP_I1;
    input CT_CAP_I2;
    input CT_CAP_I3;
    input CT_CAP_I4;
    input CT_RESN_I1;
    input CT_RESN_I2;
    input CT_RESN_I3;
    input CT_RESN_I4;
    input CT_RESP_I1;
    input CT_RESP_I2;
    input CT_RESP_I3;
    input CT_RESP_I4;
    inout [9:0] LINK_RX0;
    inout [9:0] LINK_RX1;
    inout [9:0] LINK_RX2;
    inout [9:0] LINK_RX3;
    inout [9:0] LINK_RX4;
    inout [9:0] LINK_RX5;
    inout [19:0] LINK_TX0;
    inout [19:0] LINK_TX1;
    inout [19:0] LINK_TX2;
    inout [19:0] LINK_TX3;
    inout [19:0] LINK_TX4;
    inout [19:0] LINK_TX5;
    input LOCK_E_I;
    output LOCK_O;
    input MAIN_EN_I1;
    input MAIN_EN_I2;
    input MAIN_EN_I3;
    input MAIN_EN_I4;
    input MAIN_EN_I5;
    input MAIN_EN_I6;
    input MAIN_SG_I;
    input MARG_ISV_I1;
    input MARG_ISV_I2;
    input MARG_ISV_I3;
    input MARG_ISV_I4;
    input MARG_ISV_I5;
    input MARG_IS_I1;
    input MARG_IS_I2;
    input MARG_IS_I3;
    input MARG_IS_I4;
    input MARG_SV_I1;
    input MARG_SV_I2;
    input MARG_SV_I3;
    input MARG_SV_I4;
    input MARG_SV_I5;
    input MARG_S_I1;
    input MARG_S_I2;
    input MARG_S_I3;
    input MARG_S_I4;
    input M_EYE_I;
    input OVS_E_I;
    input PLL_RN_I;
    input POST_EN_I1;
    input POST_EN_I2;
    input POST_EN_I3;
    input POST_EN_I4;
    input POST_EN_I5;
    input POST_ISV_I1;
    input POST_ISV_I2;
    input POST_ISV_I3;
    input POST_ISV_I4;
    input POST_IS_I1;
    input POST_IS_I2;
    input POST_IS_I3;
    input POST_IS_I4;
    input POST_SG_I;
    input PRE_EN_I;
    input PRE_IS_I1;
    input PRE_IS_I2;
    input PRE_IS_I3;
    input PRE_IS_I4;
    input PRE_SG_I;
    input RST_N_I;
    input RX_SEL_I1;
    input RX_SEL_I2;
    input RX_SEL_I3;
    input RX_SEL_I4;
    input RX_SEL_I5;
    input RX_SEL_I6;
    input TST_I1;
    input TST_I2;
    input TST_I3;
    input TST_I4;
    input TST_I5;
    input TST_I6;
    input TST_I7;
    input TST_I8;
    output TST_O1;
    output TST_O2;
    output TST_O3;
    output TST_O4;
    output TST_O5;
    output TST_O6;
    output TST_O7;
    output TST_O8;
    input TX_SEL_I1;
    input TX_SEL_I2;
    input TX_SEL_I3;
    input TX_SEL_I4;
    input TX_SEL_I5;
    input TX_SEL_I6;
    parameter location = "";
    parameter main_clk_to_fabric_div_en = 1'b0;
    parameter main_clk_to_fabric_div_mode = 1'b0;
    parameter main_clk_to_fabric_sel = 1'b0;
    parameter main_test = 8'b00000000;
    parameter main_use_only_usr_clock = 1'b0;
    parameter main_use_pcs_clk_2 = 1'b0;
    parameter pcs_ovs_mode = 1'b0;
    parameter pcs_pll_lock_count = 3'b000;
    parameter pcs_word_len = 2'b00;
    parameter pll_pma_cpump_n = 3'b000;
    parameter pll_pma_divf = 2'b00;
    parameter pll_pma_divf_en_n = 1'b0;
    parameter pll_pma_divm = 2'b00;
    parameter pll_pma_divm_en_n = 1'b0;
    parameter pll_pma_divn = 1'b0;
    parameter pll_pma_divn_en_n = 1'b0;
    parameter pll_pma_int_data_len = 1'b0;
    parameter pll_pma_lvds_mux = 1'b0;
    parameter pll_pma_mux_ckref = 1'b0;
    parameter rx_pma_half_step = 1'b0;
endmodule

(* blackbox *)
module NX_PMA_U(CLK_TX_I, CLK_RX_I, CLK_REF_I, DC_E_I, DC_LCSN_I1, DC_LCSN_I2, DC_LCSN_I3, DC_LCSN_I4, DC_CCSN_I, DC_WE_N_I, DC_ADD_I1, DC_ADD_I2, DC_ADD_I3, DC_ADD_I4, DC_WDATAS_I, DC_WDATA_I1, DC_WDATA_I2, DC_WDATA_I3, DC_WDATA_I4, DC_WDATA_I5, DC_WDATA_I6
, DC_WDATA_I7, DC_WDATA_I8, DC_WDATA_I9, DC_WDATA_I10, DC_WDATA_I11, DC_WDATA_I12, PLL_RN_I, PWDN_N_I, RST_N_I, DBG_S_I1, DBG_S_I2, DBG_A_I, SE_I, SCAN_I1, SCAN_I2, SCAN_I3, SCAN_I4, SCAN_I5, SCAN_I6, SCAN_I7, SCAN_I8
, CLK_O, CLK_RX_O, LOCK_O, LOCKA_O, FB_LOCK_O, CAL_OUT_O, DBG_R_O, LL_O1, LL_O2, LL_O3, LL_O4, LL_O5, LL_O6, LL_O7, LL_O8, LL_O9, LL_O10, LL_O11, LL_O12, LL_O13, LL_O14
, LL_O15, LL_O16, LL_O17, LL_O18, LL_O19, LL_O20, SCAN_O1, SCAN_O2, SCAN_O3, SCAN_O4, SCAN_O5, SCAN_O6, SCAN_O7, SCAN_O8, LINK_TX1, LINK_TX2, LINK_TX3, LINK_RX0, LINK_RX1, LINK_RX2, LINK_RX3
, LINK_TX0);
    output CAL_OUT_O;
    output CLK_O;
    input CLK_REF_I;
    input CLK_RX_I;
    output CLK_RX_O;
    input CLK_TX_I;
    input DBG_A_I;
    output DBG_R_O;
    input DBG_S_I1;
    input DBG_S_I2;
    input DC_ADD_I1;
    input DC_ADD_I2;
    input DC_ADD_I3;
    input DC_ADD_I4;
    input DC_CCSN_I;
    input DC_E_I;
    input DC_LCSN_I1;
    input DC_LCSN_I2;
    input DC_LCSN_I3;
    input DC_LCSN_I4;
    input DC_WDATAS_I;
    input DC_WDATA_I1;
    input DC_WDATA_I10;
    input DC_WDATA_I11;
    input DC_WDATA_I12;
    input DC_WDATA_I2;
    input DC_WDATA_I3;
    input DC_WDATA_I4;
    input DC_WDATA_I5;
    input DC_WDATA_I6;
    input DC_WDATA_I7;
    input DC_WDATA_I8;
    input DC_WDATA_I9;
    input DC_WE_N_I;
    output FB_LOCK_O;
    inout [9:0] LINK_RX0;
    inout [9:0] LINK_RX1;
    inout [9:0] LINK_RX2;
    inout [9:0] LINK_RX3;
    inout [19:0] LINK_TX0;
    inout [19:0] LINK_TX1;
    inout [19:0] LINK_TX2;
    inout [19:0] LINK_TX3;
    output LL_O1;
    output LL_O10;
    output LL_O11;
    output LL_O12;
    output LL_O13;
    output LL_O14;
    output LL_O15;
    output LL_O16;
    output LL_O17;
    output LL_O18;
    output LL_O19;
    output LL_O2;
    output LL_O20;
    output LL_O3;
    output LL_O4;
    output LL_O5;
    output LL_O6;
    output LL_O7;
    output LL_O8;
    output LL_O9;
    output LOCKA_O;
    output LOCK_O;
    input PLL_RN_I;
    input PWDN_N_I;
    input RST_N_I;
    input SCAN_I1;
    input SCAN_I2;
    input SCAN_I3;
    input SCAN_I4;
    input SCAN_I5;
    input SCAN_I6;
    input SCAN_I7;
    input SCAN_I8;
    output SCAN_O1;
    output SCAN_O2;
    output SCAN_O3;
    output SCAN_O4;
    output SCAN_O5;
    output SCAN_O6;
    output SCAN_O7;
    output SCAN_O8;
    input SE_I;
    parameter dyn_all_rx_pma_m_eye = 1'b0;
    parameter dyn_all_rx_pma_m_eye_coarse_ena = 1'b0;
    parameter dyn_all_rx_pma_m_eye_dn = 1'b0;
    parameter dyn_all_rx_pma_m_eye_fine_ena = 1'b0;
    parameter dyn_all_rx_pma_m_eye_step = 4'b0000;
    parameter dyn_all_rx_pma_m_eye_up = 1'b0;
    parameter dyn_all_rx_pma_threshold_1 = 5'b00000;
    parameter dyn_all_rx_pma_threshold_2 = 5'b00000;
    parameter dyn_all_rx_pma_trim_locked = 3'b000;
    parameter dyn_all_rx_pma_trim_mode = 2'b00;
    parameter dyn_all_rx_pma_trim_unlocked = 3'b000;
    parameter dyn_rx0_pma_ctle_cap_p = 4'b0000;
    parameter dyn_rx0_pma_ctle_res_p = 4'b0000;
    parameter dyn_rx0_pma_dfe_idac_tap1_n = 6'b000000;
    parameter dyn_rx0_pma_dfe_idac_tap2_n = 6'b000000;
    parameter dyn_rx0_pma_dfe_idac_tap3_n = 6'b000000;
    parameter dyn_rx0_pma_dfe_idac_tap4_n = 6'b000000;
    parameter dyn_rx0_pma_termination_cmd = 6'b000000;
    parameter dyn_rx1_pma_ctle_cap_p = 4'b0000;
    parameter dyn_rx1_pma_ctle_res_p = 4'b0000;
    parameter dyn_rx1_pma_dfe_idac_tap1_n = 6'b000000;
    parameter dyn_rx1_pma_dfe_idac_tap2_n = 6'b000000;
    parameter dyn_rx1_pma_dfe_idac_tap3_n = 6'b000000;
    parameter dyn_rx1_pma_dfe_idac_tap4_n = 6'b000000;
    parameter dyn_rx1_pma_termination_cmd = 6'b000000;
    parameter dyn_rx2_pma_ctle_cap_p = 4'b0000;
    parameter dyn_rx2_pma_ctle_res_p = 4'b0000;
    parameter dyn_rx2_pma_dfe_idac_tap1_n = 6'b000000;
    parameter dyn_rx2_pma_dfe_idac_tap2_n = 6'b000000;
    parameter dyn_rx2_pma_dfe_idac_tap3_n = 6'b000000;
    parameter dyn_rx2_pma_dfe_idac_tap4_n = 6'b000000;
    parameter dyn_rx2_pma_termination_cmd = 6'b000000;
    parameter dyn_rx3_pma_ctle_cap_p = 4'b0000;
    parameter dyn_rx3_pma_ctle_res_p = 4'b0000;
    parameter dyn_rx3_pma_dfe_idac_tap1_n = 6'b000000;
    parameter dyn_rx3_pma_dfe_idac_tap2_n = 6'b000000;
    parameter dyn_rx3_pma_dfe_idac_tap3_n = 6'b000000;
    parameter dyn_rx3_pma_dfe_idac_tap4_n = 6'b000000;
    parameter dyn_rx3_pma_termination_cmd = 6'b000000;
    parameter dyn_tx0_pma_main_en = 6'b000000;
    parameter dyn_tx0_pma_main_sign = 1'b0;
    parameter dyn_tx0_pma_margin_input = 9'b000000000;
    parameter dyn_tx0_pma_margin_sel = 9'b000000000;
    parameter dyn_tx0_pma_post_en = 5'b00000;
    parameter dyn_tx0_pma_post_sel = 8'b00000000;
    parameter dyn_tx0_pma_post_sign = 1'b0;
    parameter dyn_tx0_pma_pre_en = 1'b0;
    parameter dyn_tx0_pma_pre_sel = 4'b0000;
    parameter dyn_tx0_pma_pre_sign = 1'b0;
    parameter dyn_tx1_pma_main_en = 6'b000000;
    parameter dyn_tx1_pma_main_sign = 1'b0;
    parameter dyn_tx1_pma_margin_input = 9'b000000000;
    parameter dyn_tx1_pma_margin_sel = 9'b000000000;
    parameter dyn_tx1_pma_post_en = 5'b00000;
    parameter dyn_tx1_pma_post_sel = 8'b00000000;
    parameter dyn_tx1_pma_post_sign = 1'b0;
    parameter dyn_tx1_pma_pre_en = 1'b0;
    parameter dyn_tx1_pma_pre_sel = 4'b0000;
    parameter dyn_tx1_pma_pre_sign = 1'b0;
    parameter dyn_tx2_pma_main_en = 6'b000000;
    parameter dyn_tx2_pma_main_sign = 1'b0;
    parameter dyn_tx2_pma_margin_input = 9'b000000000;
    parameter dyn_tx2_pma_margin_sel = 9'b000000000;
    parameter dyn_tx2_pma_post_en = 5'b00000;
    parameter dyn_tx2_pma_post_sel = 8'b00000000;
    parameter dyn_tx2_pma_post_sign = 1'b0;
    parameter dyn_tx2_pma_pre_en = 1'b0;
    parameter dyn_tx2_pma_pre_sel = 4'b0000;
    parameter dyn_tx2_pma_pre_sign = 1'b0;
    parameter dyn_tx3_pma_main_en = 6'b000000;
    parameter dyn_tx3_pma_main_sign = 1'b0;
    parameter dyn_tx3_pma_margin_input = 9'b000000000;
    parameter dyn_tx3_pma_margin_sel = 9'b000000000;
    parameter dyn_tx3_pma_post_en = 5'b00000;
    parameter dyn_tx3_pma_post_sel = 8'b00000000;
    parameter dyn_tx3_pma_post_sign = 1'b0;
    parameter dyn_tx3_pma_pre_en = 1'b0;
    parameter dyn_tx3_pma_pre_sel = 4'b0000;
    parameter dyn_tx3_pma_pre_sign = 1'b0;
    parameter location = "";
    parameter main_clk_to_fabric_div_en = 1'b0;
    parameter main_clk_to_fabric_div_mode = 1'b0;
    parameter main_clk_to_fabric_sel = 1'b0;
    parameter main_rclk_to_fabric_sel = 2'b00;
    parameter main_use_only_usr_clock = 1'b0;
    parameter pcs_ovs_en = 1'b0;
    parameter pcs_ovs_mode = 1'b0;
    parameter pcs_pll_lock_ppm = 3'b000;
    parameter pcs_word_len = 2'b00;
    parameter pll_pma_ckref_ext = 1'b0;
    parameter pll_pma_cpump = 4'b0000;
    parameter pll_pma_divl = 2'b00;
    parameter pll_pma_divm = 1'b0;
    parameter pll_pma_divn = 2'b00;
    parameter pll_pma_gbx_en = 1'b0;
    parameter pll_pma_int_data_len = 1'b0;
    parameter pll_pma_lvds_en = 1'b0;
    parameter pll_pma_lvds_mux = 1'b0;
    parameter pll_pma_mux_ckref = 1'b0;
    parameter rx_usrclk_use_pcs_clk_2 = 1'b0;
    parameter test_mode = 2'b00;
    parameter tx_usrclk_use_pcs_clk_2 = 1'b0;
endmodule

(* blackbox *)
module NX_RAM(ACK, ACKC, ACKD, ACKR, BCK, BCKC, BCKD, BCKR, AI1, AI2, AI3, AI4, AI5, AI6, AI7, AI8, AI9, AI10, AI11, AI12, AI13
, AI14, AI15, AI16, AI17, AI18, AI19, AI20, AI21, AI22, AI23, AI24, BI1, BI2, BI3, BI4, BI5, BI6, BI7, BI8, BI9, BI10
, BI11, BI12, BI13, BI14, BI15, BI16, BI17, BI18, BI19, BI20, BI21, BI22, BI23, BI24, ACOR, AERR, BCOR, BERR, AO1, AO2, AO3
, AO4, AO5, AO6, AO7, AO8, AO9, AO10, AO11, AO12, AO13, AO14, AO15, AO16, AO17, AO18, AO19, AO20, AO21, AO22, AO23, AO24
, BO1, BO2, BO3, BO4, BO5, BO6, BO7, BO8, BO9, BO10, BO11, BO12, BO13, BO14, BO15, BO16, BO17, BO18, BO19, BO20, BO21
, BO22, BO23, BO24, AA1, AA2, AA3, AA4, AA5, AA6, AA7, AA8, AA9, AA10, AA11, AA12, AA13, AA14, AA15, AA16, ACS, AWE
, AR, BA1, BA2, BA3, BA4, BA5, BA6, BA7, BA8, BA9, BA10, BA11, BA12, BA13, BA14, BA15, BA16, BCS, BWE, BR);
    input AA1;
    input AA10;
    input AA11;
    input AA12;
    input AA13;
    input AA14;
    input AA15;
    input AA16;
    input AA2;
    input AA3;
    input AA4;
    input AA5;
    input AA6;
    input AA7;
    input AA8;
    input AA9;
    input ACK;
    input ACKC;
    input ACKD;
    input ACKR;
    output ACOR;
    input ACS;
    output AERR;
    input AI1;
    input AI10;
    input AI11;
    input AI12;
    input AI13;
    input AI14;
    input AI15;
    input AI16;
    input AI17;
    input AI18;
    input AI19;
    input AI2;
    input AI20;
    input AI21;
    input AI22;
    input AI23;
    input AI24;
    input AI3;
    input AI4;
    input AI5;
    input AI6;
    input AI7;
    input AI8;
    input AI9;
    output AO1;
    output AO10;
    output AO11;
    output AO12;
    output AO13;
    output AO14;
    output AO15;
    output AO16;
    output AO17;
    output AO18;
    output AO19;
    output AO2;
    output AO20;
    output AO21;
    output AO22;
    output AO23;
    output AO24;
    output AO3;
    output AO4;
    output AO5;
    output AO6;
    output AO7;
    output AO8;
    output AO9;
    input AR;
    input AWE;
    input BA1;
    input BA10;
    input BA11;
    input BA12;
    input BA13;
    input BA14;
    input BA15;
    input BA16;
    input BA2;
    input BA3;
    input BA4;
    input BA5;
    input BA6;
    input BA7;
    input BA8;
    input BA9;
    input BCK;
    input BCKC;
    input BCKD;
    input BCKR;
    output BCOR;
    input BCS;
    output BERR;
    input BI1;
    input BI10;
    input BI11;
    input BI12;
    input BI13;
    input BI14;
    input BI15;
    input BI16;
    input BI17;
    input BI18;
    input BI19;
    input BI2;
    input BI20;
    input BI21;
    input BI22;
    input BI23;
    input BI24;
    input BI3;
    input BI4;
    input BI5;
    input BI6;
    input BI7;
    input BI8;
    input BI9;
    output BO1;
    output BO10;
    output BO11;
    output BO12;
    output BO13;
    output BO14;
    output BO15;
    output BO16;
    output BO17;
    output BO18;
    output BO19;
    output BO2;
    output BO20;
    output BO21;
    output BO22;
    output BO23;
    output BO24;
    output BO3;
    output BO4;
    output BO5;
    output BO6;
    output BO7;
    output BO8;
    output BO9;
    input BR;
    input BWE;
    parameter mcka_edge = 1'b0;
    parameter mckb_edge = 1'b0;
    parameter mem_ctxt = "";
    parameter pcka_edge = 1'b0;
    parameter pckb_edge = 1'b0;
    parameter pipe_ia = 1'b0;
    parameter pipe_ib = 1'b0;
    parameter pipe_oa = 1'b0;
    parameter pipe_ob = 1'b0;
    parameter raw_config0 = 4'b0000;
    parameter raw_config1 = 16'b0000000000000000;
    parameter raw_l_enable = 1'b0;
    parameter raw_l_extend = 4'b0000;
    parameter raw_u_enable = 1'b0;
    parameter raw_u_extend = 8'b00000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_RAM_SLOWECC_1K_36_1r1w(ACK, BCK, ACOR, AERR, ACS, AWE, AR, BCS, BWE, BR, AO, AI, AA);
    input [9:0] AA;
    input ACK;
    output ACOR;
    input ACS;
    output AERR;
    input [35:0] AI;
    output [35:0] AO;
    input AR;
    input AWE;
    input BCK;
    input BCS;
    input BR;
    input BWE;
    parameter mem_ctxt = "";
endmodule

(* blackbox *)
module NX_RAM_WRAP(ACK, ACKD, ACKR, BCK, BCKD, BCKR, ACOR, AERR, BCOR, BERR, ACS, AWE, AR, BCS, BWE, BR, BI, AO, BO, AI, AA
, BA);
    input [15:0] AA;
    input ACK;
    input ACKD;
    input ACKR;
    output ACOR;
    input ACS;
    output AERR;
    input [23:0] AI;
    output [23:0] AO;
    input AR;
    input AWE;
    input [15:0] BA;
    input BCK;
    input BCKD;
    input BCKR;
    output BCOR;
    input BCS;
    output BERR;
    input [23:0] BI;
    output [23:0] BO;
    input BR;
    input BWE;
    parameter mcka_edge = 1'b0;
    parameter mckb_edge = 1'b0;
    parameter mem_ctxt = "";
    parameter pcka_edge = 1'b0;
    parameter pckb_edge = 1'b0;
    parameter pipe_ia = 1'b0;
    parameter pipe_ib = 1'b0;
    parameter pipe_oa = 1'b0;
    parameter pipe_ob = 1'b0;
    parameter raw_config0 = 4'b0000;
    parameter raw_config1 = 16'b0000000000000000;
    parameter raw_l_enable = 1'b0;
    parameter raw_l_extend = 4'b0000;
    parameter raw_u_enable = 1'b0;
    parameter raw_u_extend = 8'b00000000;
    parameter std_mode = "";
endmodule

(* blackbox *)
module NX_RB(CK1, CK2, CK3, CK4, EI1, EI2, EI3, EI4, EI5, EI6, EI7, EI8, EI9, EI10, EI11, EI12, EI13, EI14, EI15, EI16, EI17
, EI18, EI19, EI20, EI21, EI22, EI23, EI24, EI25, EI26, EI27, EI28, EI29, EI30, EI31, EI32, EI33, EI34, EI35, EI36, EI37, EI38
, EI39, EI40, EI41, EI42, EI43, EI44, EI45, EI46, EI47, EI48, EI49, EI50, EI51, EI52, EI53, EI54, EI55, EI56, EI57, EI58, EI59
, EI60, EI61, EI62, EI63, EI64, EI65, EI66, EI67, EI68, EI69, EI70, EI71, EI72, EI73, EI74, EI75, EI76, EI77, EI78, EI79, EI80
, EI81, EI82, EI83, EI84, EI85, EI86, EI87, EI88, EI89, EI90, EI91, EI92, EI93, EI94, EI95, EI96, EI97, EI98, EI99, EI100, EI101
, EI102, EI103, EI104, EI105, EI106, EI107, EI108, EI109, EI110, EI111, EI112, EI113, EI114, EI115, EI116, EI117, EI118, EI119, EI120, EI121, EI122
, EI123, EI124, EI125, EI126, EI127, EI128, EI129, EI130, EI131, EI132, EI133, EI134, EI135, EI136, EI137, EI138, EI139, EI140, EI141, EI142, EI143
, EI144, EI145, EI146, EI147, EI148, EI149, EI150, EI151, EI152, EI153, EI154, EI155, EI156, EI157, EI158, EI159, EI160, EI161, EI162, EI163, EI164
, EI165, EI166, EI167, EI168, EI169, EI170, EI171, EI172, EI173, EI174, EI175, EI176, EI177, EI178, EI179, EI180, EI181, EI182, EI183, EI184, EI185
, EI186, EI187, EI188, EI189, EI190, EI191, EI192, EI_CK, EO_CK, EO1, EO2, EO3, EO4, EO5, EO6, EO7, EO8, EO9, EO10, EO11, EO12
, EO13, EO14, EO15, EO16, EO17, EO18, EO19, EO20, EO21, EO22, EO23, EO24, EO25, EO26, EO27, EO28, EO29, EO30, EO31, EO32, EO33
, EO34, EO35, EO36, EO37, EO38, EO39, EO40, EO41, EO42, EO43, EO44, EO45, EO46, EO47, EO48, EO49, EO50, EO51, EO52, EO53, EO54
, EO55, EO56, EO57, EO58, EO59, EO60, EO61, EO62, EO63, EO64, EO65, EO66, EO67, EO68, EO69, EO70, EO71, EO72, EO73, EO74, EO75
, EO76, EO77, EO78, EO79, EO80, EO81, EO82, EO83, EO84, EO85, EO86, EO87, EO88, EO89, EO90, EO91, EO92, EO93, EO94, EO95, EO96
, EO97, EO98, EO99, EO100, EO101, EO102, EO103, EO104, EO105, EO106, EO107, EO108, EO109, EO110, EO111, EO112, EO113, EO114, EO115, EO116, EO117
, EO118, EO119, EO120, EO121, EO122, EO123, EO124, EO125, EO126, EO127, EO128, EO129, EO130, EO131, EO132, EO133, EO134, EO135, EO136, EO137, EO138
, EO139, EO140, EO141, EO142, EO143, EO144, EO145, EO146, EO147, EO148, EO149, EO150, EO151, EO152, EO153, EO154, EO155, EO156, EO157, EO158, EO159
, EO160, EO161, EO162, EO163, EO164, EO165, EO166, EO167, EO168, EO169, EO170, EO171, EO172, EO173, EO174, EO175, EO176, EO177, EO178, EO179, EO180
, EO181, EO182, EO183, EO184, EO185, EO186, EO187, EO188, EO189, EO190, EO191, EO192, FI1, FI2, FI3, FI4, FI5, FI6, FI7, FI8, FI9
, FI10, FI11, FI12, FI13, FI14, FI15, FI16, FI17, FI18, FI19, FI20, FI21, FI22, FI23, FI24, FI25, FI26, FI27, FI28, FI29, FI30
, FI31, FI32, FI33, FI34, FI35, FI36, FI37, FI38, FI39, FI40, FI41, FI42, FI43, FI44, FI45, FI46, FI47, FI48, FI49, FI50, FI51
, FI52, FI53, FI54, FI55, FI56, FI57, FI58, FI59, FI60, FI61, FI62, FI63, FI64, FI65, FI66, FI67, FI68, FI69, FI70, FI71, FI72
, FI73, FI74, FI75, FI76, FI77, FI78, FI79, FI80, FI81, FI82, FI83, FI84, FI85, FI86, FI87, FI88, FI89, FI90, FI91, FI92, FI93
, FI94, FI95, FI96, FI97, FI98, FI99, FI100, FI101, FI102, FI103, FI104, FI105, FI106, FI107, FI108, FI109, FI110, FI111, FI112, FI113, FI114
, FI115, FI116, FI117, FI118, FI119, FI120, FI121, FI122, FI123, FI124, FI125, FI126, FI127, FI128, FI129, FI130, FI131, FI132, FI133, FI134, FI135
, FI136, FI137, FI138, FI139, FI140, FI141, FI142, FI143, FI144, FI145, FI146, FI147, FI148, FI149, FI150, FI151, FI152, FI153, FI154, FI155, FI156
, FI157, FI158, FI159, FI160, FI161, FI162, FI163, FI164, FI165, FI166, FI167, FI168, FI169, FI170, FI171, FI172, FI173, FI174, FI175, FI176, FI177
, FI178, FI179, FI180, FI181, FI182, FI183, FI184, FI185, FI186, FI187, FI188, FI189, FI190, FI191, FI192, FO1, FO2, FO3, FO4, FO5, FO6
, FO7, FO8, FO9, FO10, FO11, FO12, FO13, FO14, FO15, FO16, FO17, FO18, FO19, FO20, FO21, FO22, FO23, FO24, FO25, FO26, FO27
, FO28, FO29, FO30, FO31, FO32, FO33, FO34, FO35, FO36, FO37, FO38, FO39, FO40, FO41, FO42, FO43, FO44, FO45, FO46, FO47, FO48
, FO49, FO50, FO51, FO52, FO53, FO54, FO55, FO56, FO57, FO58, FO59, FO60, FO61, FO62, FO63, FO64, FO65, FO66, FO67, FO68, FO69
, FO70, FO71, FO72, FO73, FO74, FO75, FO76, FO77, FO78, FO79, FO80, FO81, FO82, FO83, FO84, FO85, FO86, FO87, FO88, FO89, FO90
, FO91, FO92, FO93, FO94, FO95, FO96, FO97, FO98, FO99, FO100, FO101, FO102, FO103, FO104, FO105, FO106, FO107, FO108, FO109, FO110, FO111
, FO112, FO113, FO114, FO115, FO116, FO117, FO118, FO119, FO120, FO121, FO122, FO123, FO124, FO125, FO126, FO127, FO128, FO129, FO130, FO131, FO132
, FO133, FO134, FO135, FO136, FO137, FO138, FO139, FO140, FO141, FO142, FO143, FO144, FO145, FO146, FO147, FO148, FO149, FO150, FO151, FO152, FO153
, FO154, FO155, FO156, FO157, FO158, FO159, FO160, FO161, FO162, FO163, FO164, FO165, FO166, FO167, FO168, FO169, FO170, FO171, FO172, FO173, FO174
, FO175, FO176, FO177, FO178, FO179, FO180, FO181, FO182, FO183, FO184, FO185, FO186, FO187, FO188, FO189, FO190, FO191, FO192);
    input CK1;
    input CK2;
    input CK3;
    input CK4;
    input EI1;
    input EI10;
    input EI100;
    input EI101;
    input EI102;
    input EI103;
    input EI104;
    input EI105;
    input EI106;
    input EI107;
    input EI108;
    input EI109;
    input EI11;
    input EI110;
    input EI111;
    input EI112;
    input EI113;
    input EI114;
    input EI115;
    input EI116;
    input EI117;
    input EI118;
    input EI119;
    input EI12;
    input EI120;
    input EI121;
    input EI122;
    input EI123;
    input EI124;
    input EI125;
    input EI126;
    input EI127;
    input EI128;
    input EI129;
    input EI13;
    input EI130;
    input EI131;
    input EI132;
    input EI133;
    input EI134;
    input EI135;
    input EI136;
    input EI137;
    input EI138;
    input EI139;
    input EI14;
    input EI140;
    input EI141;
    input EI142;
    input EI143;
    input EI144;
    input EI145;
    input EI146;
    input EI147;
    input EI148;
    input EI149;
    input EI15;
    input EI150;
    input EI151;
    input EI152;
    input EI153;
    input EI154;
    input EI155;
    input EI156;
    input EI157;
    input EI158;
    input EI159;
    input EI16;
    input EI160;
    input EI161;
    input EI162;
    input EI163;
    input EI164;
    input EI165;
    input EI166;
    input EI167;
    input EI168;
    input EI169;
    input EI17;
    input EI170;
    input EI171;
    input EI172;
    input EI173;
    input EI174;
    input EI175;
    input EI176;
    input EI177;
    input EI178;
    input EI179;
    input EI18;
    input EI180;
    input EI181;
    input EI182;
    input EI183;
    input EI184;
    input EI185;
    input EI186;
    input EI187;
    input EI188;
    input EI189;
    input EI19;
    input EI190;
    input EI191;
    input EI192;
    input EI2;
    input EI20;
    input EI21;
    input EI22;
    input EI23;
    input EI24;
    input EI25;
    input EI26;
    input EI27;
    input EI28;
    input EI29;
    input EI3;
    input EI30;
    input EI31;
    input EI32;
    input EI33;
    input EI34;
    input EI35;
    input EI36;
    input EI37;
    input EI38;
    input EI39;
    input EI4;
    input EI40;
    input EI41;
    input EI42;
    input EI43;
    input EI44;
    input EI45;
    input EI46;
    input EI47;
    input EI48;
    input EI49;
    input EI5;
    input EI50;
    input EI51;
    input EI52;
    input EI53;
    input EI54;
    input EI55;
    input EI56;
    input EI57;
    input EI58;
    input EI59;
    input EI6;
    input EI60;
    input EI61;
    input EI62;
    input EI63;
    input EI64;
    input EI65;
    input EI66;
    input EI67;
    input EI68;
    input EI69;
    input EI7;
    input EI70;
    input EI71;
    input EI72;
    input EI73;
    input EI74;
    input EI75;
    input EI76;
    input EI77;
    input EI78;
    input EI79;
    input EI8;
    input EI80;
    input EI81;
    input EI82;
    input EI83;
    input EI84;
    input EI85;
    input EI86;
    input EI87;
    input EI88;
    input EI89;
    input EI9;
    input EI90;
    input EI91;
    input EI92;
    input EI93;
    input EI94;
    input EI95;
    input EI96;
    input EI97;
    input EI98;
    input EI99;
    output EI_CK;
    output EO1;
    output EO10;
    output EO100;
    output EO101;
    output EO102;
    output EO103;
    output EO104;
    output EO105;
    output EO106;
    output EO107;
    output EO108;
    output EO109;
    output EO11;
    output EO110;
    output EO111;
    output EO112;
    output EO113;
    output EO114;
    output EO115;
    output EO116;
    output EO117;
    output EO118;
    output EO119;
    output EO12;
    output EO120;
    output EO121;
    output EO122;
    output EO123;
    output EO124;
    output EO125;
    output EO126;
    output EO127;
    output EO128;
    output EO129;
    output EO13;
    output EO130;
    output EO131;
    output EO132;
    output EO133;
    output EO134;
    output EO135;
    output EO136;
    output EO137;
    output EO138;
    output EO139;
    output EO14;
    output EO140;
    output EO141;
    output EO142;
    output EO143;
    output EO144;
    output EO145;
    output EO146;
    output EO147;
    output EO148;
    output EO149;
    output EO15;
    output EO150;
    output EO151;
    output EO152;
    output EO153;
    output EO154;
    output EO155;
    output EO156;
    output EO157;
    output EO158;
    output EO159;
    output EO16;
    output EO160;
    output EO161;
    output EO162;
    output EO163;
    output EO164;
    output EO165;
    output EO166;
    output EO167;
    output EO168;
    output EO169;
    output EO17;
    output EO170;
    output EO171;
    output EO172;
    output EO173;
    output EO174;
    output EO175;
    output EO176;
    output EO177;
    output EO178;
    output EO179;
    output EO18;
    output EO180;
    output EO181;
    output EO182;
    output EO183;
    output EO184;
    output EO185;
    output EO186;
    output EO187;
    output EO188;
    output EO189;
    output EO19;
    output EO190;
    output EO191;
    output EO192;
    output EO2;
    output EO20;
    output EO21;
    output EO22;
    output EO23;
    output EO24;
    output EO25;
    output EO26;
    output EO27;
    output EO28;
    output EO29;
    output EO3;
    output EO30;
    output EO31;
    output EO32;
    output EO33;
    output EO34;
    output EO35;
    output EO36;
    output EO37;
    output EO38;
    output EO39;
    output EO4;
    output EO40;
    output EO41;
    output EO42;
    output EO43;
    output EO44;
    output EO45;
    output EO46;
    output EO47;
    output EO48;
    output EO49;
    output EO5;
    output EO50;
    output EO51;
    output EO52;
    output EO53;
    output EO54;
    output EO55;
    output EO56;
    output EO57;
    output EO58;
    output EO59;
    output EO6;
    output EO60;
    output EO61;
    output EO62;
    output EO63;
    output EO64;
    output EO65;
    output EO66;
    output EO67;
    output EO68;
    output EO69;
    output EO7;
    output EO70;
    output EO71;
    output EO72;
    output EO73;
    output EO74;
    output EO75;
    output EO76;
    output EO77;
    output EO78;
    output EO79;
    output EO8;
    output EO80;
    output EO81;
    output EO82;
    output EO83;
    output EO84;
    output EO85;
    output EO86;
    output EO87;
    output EO88;
    output EO89;
    output EO9;
    output EO90;
    output EO91;
    output EO92;
    output EO93;
    output EO94;
    output EO95;
    output EO96;
    output EO97;
    output EO98;
    output EO99;
    output EO_CK;
    input FI1;
    input FI10;
    input FI100;
    input FI101;
    input FI102;
    input FI103;
    input FI104;
    input FI105;
    input FI106;
    input FI107;
    input FI108;
    input FI109;
    input FI11;
    input FI110;
    input FI111;
    input FI112;
    input FI113;
    input FI114;
    input FI115;
    input FI116;
    input FI117;
    input FI118;
    input FI119;
    input FI12;
    input FI120;
    input FI121;
    input FI122;
    input FI123;
    input FI124;
    input FI125;
    input FI126;
    input FI127;
    input FI128;
    input FI129;
    input FI13;
    input FI130;
    input FI131;
    input FI132;
    input FI133;
    input FI134;
    input FI135;
    input FI136;
    input FI137;
    input FI138;
    input FI139;
    input FI14;
    input FI140;
    input FI141;
    input FI142;
    input FI143;
    input FI144;
    input FI145;
    input FI146;
    input FI147;
    input FI148;
    input FI149;
    input FI15;
    input FI150;
    input FI151;
    input FI152;
    input FI153;
    input FI154;
    input FI155;
    input FI156;
    input FI157;
    input FI158;
    input FI159;
    input FI16;
    input FI160;
    input FI161;
    input FI162;
    input FI163;
    input FI164;
    input FI165;
    input FI166;
    input FI167;
    input FI168;
    input FI169;
    input FI17;
    input FI170;
    input FI171;
    input FI172;
    input FI173;
    input FI174;
    input FI175;
    input FI176;
    input FI177;
    input FI178;
    input FI179;
    input FI18;
    input FI180;
    input FI181;
    input FI182;
    input FI183;
    input FI184;
    input FI185;
    input FI186;
    input FI187;
    input FI188;
    input FI189;
    input FI19;
    input FI190;
    input FI191;
    input FI192;
    input FI2;
    input FI20;
    input FI21;
    input FI22;
    input FI23;
    input FI24;
    input FI25;
    input FI26;
    input FI27;
    input FI28;
    input FI29;
    input FI3;
    input FI30;
    input FI31;
    input FI32;
    input FI33;
    input FI34;
    input FI35;
    input FI36;
    input FI37;
    input FI38;
    input FI39;
    input FI4;
    input FI40;
    input FI41;
    input FI42;
    input FI43;
    input FI44;
    input FI45;
    input FI46;
    input FI47;
    input FI48;
    input FI49;
    input FI5;
    input FI50;
    input FI51;
    input FI52;
    input FI53;
    input FI54;
    input FI55;
    input FI56;
    input FI57;
    input FI58;
    input FI59;
    input FI6;
    input FI60;
    input FI61;
    input FI62;
    input FI63;
    input FI64;
    input FI65;
    input FI66;
    input FI67;
    input FI68;
    input FI69;
    input FI7;
    input FI70;
    input FI71;
    input FI72;
    input FI73;
    input FI74;
    input FI75;
    input FI76;
    input FI77;
    input FI78;
    input FI79;
    input FI8;
    input FI80;
    input FI81;
    input FI82;
    input FI83;
    input FI84;
    input FI85;
    input FI86;
    input FI87;
    input FI88;
    input FI89;
    input FI9;
    input FI90;
    input FI91;
    input FI92;
    input FI93;
    input FI94;
    input FI95;
    input FI96;
    input FI97;
    input FI98;
    input FI99;
    output FO1;
    output FO10;
    output FO100;
    output FO101;
    output FO102;
    output FO103;
    output FO104;
    output FO105;
    output FO106;
    output FO107;
    output FO108;
    output FO109;
    output FO11;
    output FO110;
    output FO111;
    output FO112;
    output FO113;
    output FO114;
    output FO115;
    output FO116;
    output FO117;
    output FO118;
    output FO119;
    output FO12;
    output FO120;
    output FO121;
    output FO122;
    output FO123;
    output FO124;
    output FO125;
    output FO126;
    output FO127;
    output FO128;
    output FO129;
    output FO13;
    output FO130;
    output FO131;
    output FO132;
    output FO133;
    output FO134;
    output FO135;
    output FO136;
    output FO137;
    output FO138;
    output FO139;
    output FO14;
    output FO140;
    output FO141;
    output FO142;
    output FO143;
    output FO144;
    output FO145;
    output FO146;
    output FO147;
    output FO148;
    output FO149;
    output FO15;
    output FO150;
    output FO151;
    output FO152;
    output FO153;
    output FO154;
    output FO155;
    output FO156;
    output FO157;
    output FO158;
    output FO159;
    output FO16;
    output FO160;
    output FO161;
    output FO162;
    output FO163;
    output FO164;
    output FO165;
    output FO166;
    output FO167;
    output FO168;
    output FO169;
    output FO17;
    output FO170;
    output FO171;
    output FO172;
    output FO173;
    output FO174;
    output FO175;
    output FO176;
    output FO177;
    output FO178;
    output FO179;
    output FO18;
    output FO180;
    output FO181;
    output FO182;
    output FO183;
    output FO184;
    output FO185;
    output FO186;
    output FO187;
    output FO188;
    output FO189;
    output FO19;
    output FO190;
    output FO191;
    output FO192;
    output FO2;
    output FO20;
    output FO21;
    output FO22;
    output FO23;
    output FO24;
    output FO25;
    output FO26;
    output FO27;
    output FO28;
    output FO29;
    output FO3;
    output FO30;
    output FO31;
    output FO32;
    output FO33;
    output FO34;
    output FO35;
    output FO36;
    output FO37;
    output FO38;
    output FO39;
    output FO4;
    output FO40;
    output FO41;
    output FO42;
    output FO43;
    output FO44;
    output FO45;
    output FO46;
    output FO47;
    output FO48;
    output FO49;
    output FO5;
    output FO50;
    output FO51;
    output FO52;
    output FO53;
    output FO54;
    output FO55;
    output FO56;
    output FO57;
    output FO58;
    output FO59;
    output FO6;
    output FO60;
    output FO61;
    output FO62;
    output FO63;
    output FO64;
    output FO65;
    output FO66;
    output FO67;
    output FO68;
    output FO69;
    output FO7;
    output FO70;
    output FO71;
    output FO72;
    output FO73;
    output FO74;
    output FO75;
    output FO76;
    output FO77;
    output FO78;
    output FO79;
    output FO8;
    output FO80;
    output FO81;
    output FO82;
    output FO83;
    output FO84;
    output FO85;
    output FO86;
    output FO87;
    output FO88;
    output FO89;
    output FO9;
    output FO90;
    output FO91;
    output FO92;
    output FO93;
    output FO94;
    output FO95;
    output FO96;
    output FO97;
    output FO98;
    output FO99;
    parameter inputBypass = 24'b000000000000000000000000;
    parameter inputClk = 2'b00;
    parameter inputContext = "";
    parameter outputBypass = 24'b000000000000000000000000;
    parameter outputClk = 2'b00;
    parameter outputContext = "";
endmodule

(* blackbox *)
module NX_RB_WRAP(EI_CK, EO_CK, CK, EO, EI, FI, FO);
    input [3:0] CK;
    input [191:0] EI;
    output EI_CK;
    output [191:0] EO;
    output EO_CK;
    input [191:0] FI;
    output [191:0] FO;
    parameter inputBypass = 24'b000000000000000000000000;
    parameter inputClk = 2'b00;
    parameter inputContext = "";
    parameter outputBypass = 24'b000000000000000000000000;
    parameter outputClk = 2'b00;
    parameter outputContext = "";
endmodule

(* blackbox *)
module NX_RFB(RCK, WCK, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, COR, ERR, O1
, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, RA1, RA2, RA3, RA4, RA5, RA6
, RE, WA1, WA2, WA3, WA4, WA5, WA6, WE);
    output COR;
    output ERR;
    input I1;
    input I10;
    input I11;
    input I12;
    input I13;
    input I14;
    input I15;
    input I16;
    input I2;
    input I3;
    input I4;
    input I5;
    input I6;
    input I7;
    input I8;
    input I9;
    output O1;
    output O10;
    output O11;
    output O12;
    output O13;
    output O14;
    output O15;
    output O16;
    output O2;
    output O3;
    output O4;
    output O5;
    output O6;
    output O7;
    output O8;
    output O9;
    input RA1;
    input RA2;
    input RA3;
    input RA4;
    input RA5;
    input RA6;
    input RCK;
    input RE;
    input WA1;
    input WA2;
    input WA3;
    input WA4;
    input WA5;
    input WA6;
    input WCK;
    input WE;
    parameter addr_mask = 5'b00000;
    parameter mem_ctxt = "";
    parameter rck_edge = 1'b0;
    parameter wck_edge = 1'b0;
    parameter we_mask = 1'b0;
    parameter wea_mask = 1'b0;
endmodule

(* blackbox *)
module NX_RFBDP_U_WRAP(WCK, WE, WEA, I, O, RA, WA);
    input [17:0] I;
    output [17:0] O;
    input [4:0] RA;
    input [4:0] WA;
    input WCK;
    input WE;
    input WEA;
    parameter mem_ctxt = "";
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_RFBSP_U_WRAP(WCK, WE, WEA, I, O, WA);
    input [17:0] I;
    output [17:0] O;
    input [4:0] WA;
    input WCK;
    input WE;
    input WEA;
    parameter mem_ctxt = "";
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_RFB_L(RCK, WCK, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, COR, ERR, O1
, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, RA1, RA2, RA3, RA4, RA5, RA6
, RE, WA1, WA2, WA3, WA4, WA5, WA6, WE);
    output COR;
    output ERR;
    input I1;
    input I10;
    input I11;
    input I12;
    input I13;
    input I14;
    input I15;
    input I16;
    input I2;
    input I3;
    input I4;
    input I5;
    input I6;
    input I7;
    input I8;
    input I9;
    output O1;
    output O10;
    output O11;
    output O12;
    output O13;
    output O14;
    output O15;
    output O16;
    output O2;
    output O3;
    output O4;
    output O5;
    output O6;
    output O7;
    output O8;
    output O9;
    input RA1;
    input RA2;
    input RA3;
    input RA4;
    input RA5;
    input RA6;
    input RCK;
    input RE;
    input WA1;
    input WA2;
    input WA3;
    input WA4;
    input WA5;
    input WA6;
    input WCK;
    input WE;
    parameter mem_ctxt = "";
    parameter mode = 0;
    parameter rck_edge = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_RFB_L_WRAP(RCK, WCK, COR, ERR, RE, WE, I, O, RA, WA);
    output COR;
    output ERR;
    input [15:0] I;
    output [15:0] O;
    input [5:0] RA;
    input RCK;
    input RE;
    input [5:0] WA;
    input WCK;
    input WE;
    parameter mem_ctxt = "";
    parameter mode = 0;
    parameter rck_edge = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_RFB_M(RCK, WCK, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, COR, ERR, O1
, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, RA1, RA2, RA3, RA4, RA5, RA6
, RE, WA1, WA2, WA3, WA4, WA5, WA6, WE);
    output COR;
    output ERR;
    input I1;
    input I10;
    input I11;
    input I12;
    input I13;
    input I14;
    input I15;
    input I16;
    input I2;
    input I3;
    input I4;
    input I5;
    input I6;
    input I7;
    input I8;
    input I9;
    output O1;
    output O10;
    output O11;
    output O12;
    output O13;
    output O14;
    output O15;
    output O16;
    output O2;
    output O3;
    output O4;
    output O5;
    output O6;
    output O7;
    output O8;
    output O9;
    input RA1;
    input RA2;
    input RA3;
    input RA4;
    input RA5;
    input RA6;
    input RCK;
    input RE;
    input WA1;
    input WA2;
    input WA3;
    input WA4;
    input WA5;
    input WA6;
    input WCK;
    input WE;
    parameter mem_ctxt = "";
    parameter rck_edge = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_RFB_U(WCK, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20
, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, I32, I33, I34, I35, I36, O1, O2, O3, O4, O5
, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15, O16, O17, O18, O19, O20, O21, O22, O23, O24, O25, O26
, O27, O28, O29, O30, O31, O32, O33, O34, O35, O36, RA1, RA2, RA3, RA4, RA5, RA6, RA7, RA8, RA9, RA10, WA1
, WA2, WA3, WA4, WA5, WA6, WE, WEA);
    input I1;
    input I10;
    input I11;
    input I12;
    input I13;
    input I14;
    input I15;
    input I16;
    input I17;
    input I18;
    input I19;
    input I2;
    input I20;
    input I21;
    input I22;
    input I23;
    input I24;
    input I25;
    input I26;
    input I27;
    input I28;
    input I29;
    input I3;
    input I30;
    input I31;
    input I32;
    input I33;
    input I34;
    input I35;
    input I36;
    input I4;
    input I5;
    input I6;
    input I7;
    input I8;
    input I9;
    output O1;
    output O10;
    output O11;
    output O12;
    output O13;
    output O14;
    output O15;
    output O16;
    output O17;
    output O18;
    output O19;
    output O2;
    output O20;
    output O21;
    output O22;
    output O23;
    output O24;
    output O25;
    output O26;
    output O27;
    output O28;
    output O29;
    output O3;
    output O30;
    output O31;
    output O32;
    output O33;
    output O34;
    output O35;
    output O36;
    output O4;
    output O5;
    output O6;
    output O7;
    output O8;
    output O9;
    input RA1;
    input RA10;
    input RA2;
    input RA3;
    input RA4;
    input RA5;
    input RA6;
    input RA7;
    input RA8;
    input RA9;
    input WA1;
    input WA2;
    input WA3;
    input WA4;
    input WA5;
    input WA6;
    input WCK;
    input WE;
    input WEA;
    parameter mem_ctxt = "";
    parameter mode = 0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_RFB_WRAP(RCK, WCK, COR, ERR, RE, WE, I, O, RA, WA);
    output COR;
    output ERR;
    input [15:0] I;
    output [15:0] O;
    input [5:0] RA;
    input RCK;
    input RE;
    input [5:0] WA;
    input WCK;
    input WE;
    parameter mem_ctxt = "";
    parameter rck_edge = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_SER(FCK, SCK, R, IO, DCK, DRL, I, DS, DRA, DRI, DRO, DID);
    input DCK;
    output [5:0] DID;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    input FCK;
    input [4:0] I;
    output IO;
    input R;
    input SCK;
    parameter data_size = 5;
    parameter differential = "";
    parameter drive = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter slewRate = "";
    parameter spath_dynamic = 1'b0;
    parameter standard = "";
endmodule

(* blackbox *)
module NX_SERDES(FCK, SCK, RTX, RRX, CI, CCK, CL, CR, IO, DCK, DRL, DIG, FZ, FLD, FLG, I, O, DS, DRA, DRI, DRO
, DID);
    input CCK;
    input CI;
    input CL;
    input CR;
    input DCK;
    output [5:0] DID;
    input DIG;
    input [5:0] DRA;
    input [5:0] DRI;
    input DRL;
    output [5:0] DRO;
    input [1:0] DS;
    input FCK;
    output FLD;
    output FLG;
    input FZ;
    input [4:0] I;
    inout IO;
    output [4:0] O;
    input RRX;
    input RTX;
    input SCK;
    parameter cpath_registered = 1'b0;
    parameter data_size = 5;
    parameter differential = "";
    parameter dpath_dynamic = 1'b0;
    parameter drive = "";
    parameter inputDelayLine = "";
    parameter inputSignalSlope = "";
    parameter location = "";
    parameter locked = 1'b0;
    parameter outputCapacity = "";
    parameter outputDelayLine = "";
    parameter slewRate = "";
    parameter spath_dynamic = 1'b0;
    parameter standard = "";
    parameter termination = "";
    parameter terminationReference = "";
    parameter turbo = "";
    parameter weakTermination = "";
endmodule

(* blackbox *)
module NX_WFG(SI, ZI, RDY, SO, ZO);
    input RDY;
    input SI;
    output SO;
    input ZI;
    output ZO;
    parameter delay = 0;
    parameter delay_on = 1'b0;
    parameter location = "";
    parameter mode = 1'b0;
    parameter pattern = 16'b0000000000000000;
    parameter pattern_end = 1;
    parameter wfg_edge = 1'b0;
endmodule

(* blackbox *)
module NX_WFG_L(R, SI, ZI, RDY, SO, ZO);
    input R;
    input RDY;
    input SI;
    output SO;
    input ZI;
    output ZO;
    parameter delay = 0;
    parameter delay_on = 1'b0;
    parameter location = "";
    parameter mode = 1'b0;
    parameter pattern = 16'b0000000000000000;
    parameter pattern_end = 1;
    parameter wfg_edge = 1'b0;
endmodule

(* blackbox *)
module NX_WFG_U(R, SI, ZI, SO, ZO);
    input R;
    input SI;
    output SO;
    input ZI;
    output ZO;
    parameter delay = 0;
    parameter delay_on = 1'b0;
    parameter div_phase = 1'b0;
    parameter div_ratio = 0;
    parameter location = "";
    parameter mode = 0;
    parameter pattern = 16'b0000000000000000;
    parameter pattern_end = 0;
    parameter reset_on_cal_lock_n = 1'b0;
    parameter reset_on_pll_lock_n = 1'b0;
    parameter reset_on_pll_locka_n = 1'b0;
    parameter wfg_edge = 1'b0;
endmodule

(* blackbox *)
module NX_XCDC_U(CK1, CK2, ASRSTI, ADRSTI, ASRSTO, ADRSTO, BSRSTI, BDRSTI, BSRSTO, BDRSTO, CSRSTI, CDRSTI, CSRSTO, CDRSTO, DSRSTI, DDRSTI, DSRSTO, DDRSTO, BI, CI, CO
, AO, BO, AI, DI, DO);
    input ADRSTI;
    output ADRSTO;
    input [5:0] AI;
    output [5:0] AO;
    input ASRSTI;
    output ASRSTO;
    input BDRSTI;
    output BDRSTO;
    input [5:0] BI;
    output [5:0] BO;
    input BSRSTI;
    output BSRSTO;
    input CDRSTI;
    output CDRSTO;
    input [5:0] CI;
    input CK1;
    input CK2;
    output [5:0] CO;
    input CSRSTI;
    output CSRSTO;
    input DDRSTI;
    output DDRSTO;
    input [5:0] DI;
    output [5:0] DO;
    input DSRSTI;
    output DSRSTO;
    parameter ack_sel = 1'b0;
    parameter bck_sel = 1'b0;
    parameter cck_sel = 1'b0;
    parameter ck0_edge = 1'b0;
    parameter ck1_edge = 1'b0;
    parameter dck_sel = 1'b0;
    parameter link_BA = 1'b0;
    parameter link_CB = 1'b0;
    parameter link_DC = 1'b0;
    parameter use_adest_arst = 1'b0;
    parameter use_asrc_arst = 1'b0;
    parameter use_bdest_arst = 1'b0;
    parameter use_bsrc_arst = 1'b0;
    parameter use_cdest_arst = 1'b0;
    parameter use_csrc_arst = 1'b0;
    parameter use_ddest_arst = 1'b0;
    parameter use_dsrc_arst = 1'b0;
endmodule

(* blackbox *)
module NX_XFIFO_32x36(RCK, WCK, WE, WEA, WRSTI, WEQ, RRSTI, REQ, I, O, WAI, WAO, RAI, RAO);
    input [35:0] I;
    output [35:0] O;
    input [5:0] RAI;
    output [5:0] RAO;
    input RCK;
    output REQ;
    input RRSTI;
    input [5:0] WAI;
    output [5:0] WAO;
    input WCK;
    input WE;
    input WEA;
    output WEQ;
    input WRSTI;
    parameter rck_edge = 1'b0;
    parameter read_addr_inv = 7'b0000000;
    parameter use_read_arst = 1'b0;
    parameter use_write_arst = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_XFIFO_64x18(RCK, WCK, WE, WEA, WRSTI, RRSTI, I, O, WEQ, REQ, WAI, WAO, RAI, RAO);
    input [17:0] I;
    output [17:0] O;
    input [6:0] RAI;
    output [6:0] RAO;
    input RCK;
    output [1:0] REQ;
    input RRSTI;
    input [6:0] WAI;
    output [6:0] WAO;
    input WCK;
    input WE;
    input WEA;
    output [1:0] WEQ;
    input WRSTI;
    parameter rck_edge = 1'b0;
    parameter read_addr_inv = 7'b0000000;
    parameter use_read_arst = 1'b0;
    parameter use_write_arst = 1'b0;
    parameter wck_edge = 1'b0;
endmodule

(* blackbox *)
module NX_XRFB_2R_1W(WCK, WE, WEA, I, AO, BO, WA, ARA, BRA);
    output [17:0] AO;
    input [4:0] ARA;
    output [17:0] BO;
    input [4:0] BRA;
    input [17:0] I;
    input [4:0] WA;
    input WCK;
    input WE;
    input WEA;
    parameter mem_ctxt = "";
    parameter wck_edge = 1'b0;
endmodule

//(* blackbox *)
//module NX_XRFB_32x36(WCK, WE, WEA, I, O, RA, WA);
//    input [35:0] I;
//    output [35:0] O;
//    input [4:0] RA;
//    input [4:0] WA;
//    input WCK;
//    input WE;
//    input WEA;
//    parameter mem_ctxt = "";
//    parameter wck_edge = 1'b0;
//endmodule
//
//(* blackbox *)
//module NX_XRFB_64x18(WCK, WE, WEA, I, O, RA, WA);
//    input [17:0] I;
//    output [17:0] O;
//    input [5:0] RA;
//    input [5:0] WA;
//    input WCK;
//    input WE;
//    input WEA;
//    parameter mem_ctxt = "";
//    parameter wck_edge = 1'b0;
//endmodule

(* blackbox *)
module SMACC24x18_1DSP(clk, rst, A, B, Z);
    input [23:0] A;
    input [17:0] B;
    output [55:0] Z;
    input clk;
    input rst;
    parameter g_pipe = 1;
endmodule

(* blackbox *)
module SMACC24x32_2DSP(clk, rst, A, B, Z);
    input [23:0] A;
    input [31:0] B;
    output [55:0] Z;
    input clk;
    input rst;
    parameter g_pipe = 1;
endmodule

(* blackbox *)
module SMACC24x32_enable_2DSP(clk, rst, we, A, B, Z);
    input [23:0] A;
    input [31:0] B;
    output [55:0] Z;
    input clk;
    input rst;
    input we;
    parameter STAGE_1 = "false";
    parameter STAGE_2 = "false";
    parameter STAGE_3 = "false";
    parameter STAGE_4 = "false";
endmodule

(* blackbox *)
module SMUL24x32_2DSP(clk, rst, A, B, Z);
    input [23:0] A;
    input [31:0] B;
    output [54:0] Z;
    input clk;
    input rst;
    parameter g_pipe = 1;
endmodule

(* blackbox *)
module SMUL24x32_2DSP_ACC_2DSP(clk, rst, we, A, B, Z);
    input [23:0] A;
    input [31:0] B;
    output [97:0] Z;
    input clk;
    input rst;
    input we;
    parameter STAGE_1 = "false";
    parameter STAGE_2 = "false";
    parameter STAGE_3 = "false";
endmodule

(* blackbox *)
module SMUL24x32_2DSP_ACC_2DSP_L(clk, rst, we, A, B, Z);
    input [23:0] A;
    input [31:0] B;
    output [91:0] Z;
    input clk;
    input rst;
    input we;
endmodule

(* blackbox *)
module SMUL47x35_4DSP(clk, rst, A, B, Z);
    input [46:0] A;
    input [34:0] B;
    output [80:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMADD24_2DSP(clk, rst, A, B, C, Z);
    input [23:0] A;
    input [31:0] B;
    input [55:0] C;
    output [55:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMUL24x32_1DSP_2CYCLES(clk, rst, A, B, Z);
    input [23:0] A;
    input [15:0] B;
    output [55:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMUL24x32_2DSP(clk, rst, A, B, Z);
    input [23:0] A;
    input [31:0] B;
    output [55:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMUL24x36_1DSP_2CYCLES(clk, rst, A, B, Z);
    input [23:0] A;
    input [17:0] B;
    output [59:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMUL24x36_2DSP(clk, rst, A, B, Z);
    input [23:0] A;
    input [35:0] B;
    output [59:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMUL48x36_1DSP_4CYCLES(clk, rst, A, B, Z);
    input [23:0] A;
    input [17:0] B;
    output [83:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule

(* blackbox *)
module UMUL48x36_4DSP(clk, rst, A, B, Z);
    input [47:0] A;
    input [35:0] B;
    output [83:0] Z;
    input clk;
    input rst;
    parameter piped = "true";
endmodule
