// Created by cells_xtra.py from Xilinx models

module PCIE_2_0 (...);
    parameter [11:0] AER_BASE_PTR = 12'h128;
    parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [15:0] AER_CAP_ID = 16'h0001;
    parameter [4:0] AER_CAP_INT_MSG_NUM_MSI = 5'h0A;
    parameter [4:0] AER_CAP_INT_MSG_NUM_MSIX = 5'h15;
    parameter [11:0] AER_CAP_NEXTPTR = 12'h160;
    parameter AER_CAP_ON = "FALSE";
    parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
    parameter [3:0] AER_CAP_VERSION = 4'h1;
    parameter ALLOW_X8_GEN2 = "FALSE";
    parameter [31:0] BAR0 = 32'hFFFFFF00;
    parameter [31:0] BAR1 = 32'hFFFF0000;
    parameter [31:0] BAR2 = 32'hFFFF000C;
    parameter [31:0] BAR3 = 32'hFFFFFFFF;
    parameter [31:0] BAR4 = 32'h00000000;
    parameter [31:0] BAR5 = 32'h00000000;
    parameter [7:0] CAPABILITIES_PTR = 8'h40;
    parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
    parameter [23:0] CLASS_CODE = 24'h000000;
    parameter CMD_INTX_IMPLEMENTED = "TRUE";
    parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
    parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
    parameter [6:0] CRM_MODULE_RSTS = 7'h00;
    parameter [15:0] DEVICE_ID = 16'h0007;
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
    parameter integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
    parameter integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
    parameter integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
    parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
    parameter integer DEV_CAP_RSVD_14_12 = 0;
    parameter integer DEV_CAP_RSVD_17_16 = 0;
    parameter integer DEV_CAP_RSVD_31_29 = 0;
    parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
    parameter DISABLE_ASPM_L1_TIMER = "FALSE";
    parameter DISABLE_BAR_FILTERING = "FALSE";
    parameter DISABLE_ID_CHECK = "FALSE";
    parameter DISABLE_LANE_REVERSAL = "FALSE";
    parameter DISABLE_RX_TC_FILTER = "FALSE";
    parameter DISABLE_SCRAMBLING = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [11:0] DSN_BASE_PTR = 12'h100;
    parameter [15:0] DSN_CAP_ID = 16'h0003;
    parameter [11:0] DSN_CAP_NEXTPTR = 12'h000;
    parameter DSN_CAP_ON = "TRUE";
    parameter [3:0] DSN_CAP_VERSION = 4'h1;
    parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
    parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
    parameter ENTER_RVRY_EI_L0 = "TRUE";
    parameter EXIT_LOOPBACK_ON_EI = "TRUE";
    parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
    parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
    parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
    parameter [7:0] HEADER_TYPE = 8'h00;
    parameter [4:0] INFER_EI = 5'h00;
    parameter [7:0] INTERRUPT_PIN = 8'h01;
    parameter IS_SWITCH = "FALSE";
    parameter [9:0] LAST_CONFIG_DWORD = 10'h042;
    parameter integer LINK_CAP_ASPM_SUPPORT = 1;
    parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
    parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
    parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
    parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
    parameter integer LINK_CAP_RSVD_23_22 = 0;
    parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
    parameter integer LINK_CONTROL_RCB = 0;
    parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
    parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
    parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
    parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
    parameter [7:0] MSIX_BASE_PTR = 8'h9C;
    parameter [7:0] MSIX_CAP_ID = 8'h11;
    parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
    parameter MSIX_CAP_ON = "FALSE";
    parameter integer MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] MSI_BASE_PTR = 8'h48;
    parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
    parameter [7:0] MSI_CAP_ID = 8'h05;
    parameter integer MSI_CAP_MULTIMSGCAP = 0;
    parameter integer MSI_CAP_MULTIMSG_EXTENSION = 0;
    parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
    parameter MSI_CAP_ON = "FALSE";
    parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
    parameter integer N_FTS_COMCLK_GEN1 = 255;
    parameter integer N_FTS_COMCLK_GEN2 = 255;
    parameter integer N_FTS_GEN1 = 255;
    parameter integer N_FTS_GEN2 = 255;
    parameter [7:0] PCIE_BASE_PTR = 8'h60;
    parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
    parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
    parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
    parameter [4:0] PCIE_CAP_INT_MSG_NUM = 5'h00;
    parameter [7:0] PCIE_CAP_NEXTPTR = 8'h00;
    parameter PCIE_CAP_ON = "TRUE";
    parameter integer PCIE_CAP_RSVD_15_14 = 0;
    parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
    parameter integer PCIE_REVISION = 2;
    parameter integer PGL0_LANE = 0;
    parameter integer PGL1_LANE = 1;
    parameter integer PGL2_LANE = 2;
    parameter integer PGL3_LANE = 3;
    parameter integer PGL4_LANE = 4;
    parameter integer PGL5_LANE = 5;
    parameter integer PGL6_LANE = 6;
    parameter integer PGL7_LANE = 7;
    parameter integer PL_AUTO_CONFIG = 0;
    parameter PL_FAST_TRAIN = "FALSE";
    parameter [7:0] PM_BASE_PTR = 8'h40;
    parameter integer PM_CAP_AUXCURRENT = 0;
    parameter PM_CAP_D1SUPPORT = "TRUE";
    parameter PM_CAP_D2SUPPORT = "TRUE";
    parameter PM_CAP_DSI = "FALSE";
    parameter [7:0] PM_CAP_ID = 8'h01;
    parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
    parameter PM_CAP_ON = "TRUE";
    parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
    parameter PM_CAP_PME_CLOCK = "FALSE";
    parameter integer PM_CAP_RSVD_04 = 0;
    parameter integer PM_CAP_VERSION = 3;
    parameter PM_CSR_B2B3 = "FALSE";
    parameter PM_CSR_BPCCEN = "FALSE";
    parameter PM_CSR_NOSOFTRST = "TRUE";
    parameter [7:0] PM_DATA0 = 8'h01;
    parameter [7:0] PM_DATA1 = 8'h01;
    parameter [7:0] PM_DATA2 = 8'h01;
    parameter [7:0] PM_DATA3 = 8'h01;
    parameter [7:0] PM_DATA4 = 8'h01;
    parameter [7:0] PM_DATA5 = 8'h01;
    parameter [7:0] PM_DATA6 = 8'h01;
    parameter [7:0] PM_DATA7 = 8'h01;
    parameter [1:0] PM_DATA_SCALE0 = 2'h1;
    parameter [1:0] PM_DATA_SCALE1 = 2'h1;
    parameter [1:0] PM_DATA_SCALE2 = 2'h1;
    parameter [1:0] PM_DATA_SCALE3 = 2'h1;
    parameter [1:0] PM_DATA_SCALE4 = 2'h1;
    parameter [1:0] PM_DATA_SCALE5 = 2'h1;
    parameter [1:0] PM_DATA_SCALE6 = 2'h1;
    parameter [1:0] PM_DATA_SCALE7 = 2'h1;
    parameter integer RECRC_CHK = 0;
    parameter RECRC_CHK_TRIM = "FALSE";
    parameter [7:0] REVISION_ID = 8'h00;
    parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
    parameter SELECT_DLL_IF = "FALSE";
    parameter SIM_VERSION = "1.0";
    parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
    parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
    parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
    parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
    parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
    parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
    parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
    parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
    parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
    parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
    parameter integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
    parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter [15:0] SUBSYSTEM_ID = 16'h0007;
    parameter [15:0] SUBSYSTEM_VENDOR_ID = 16'h10EE;
    parameter TL_RBYPASS = "FALSE";
    parameter integer TL_RX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_RX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_RX_RAM_WRITE_LATENCY = 0;
    parameter TL_TFC_DISABLE = "FALSE";
    parameter TL_TX_CHECKS_DISABLE = "FALSE";
    parameter integer TL_TX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_TX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_TX_RAM_WRITE_LATENCY = 0;
    parameter UPCONFIG_CAPABLE = "TRUE";
    parameter UPSTREAM_FACING = "TRUE";
    parameter UR_INV_REQ = "TRUE";
    parameter integer USER_CLK_FREQ = 3;
    parameter VC0_CPL_INFINITE = "TRUE";
    parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
    parameter integer VC0_TOTAL_CREDITS_CD = 127;
    parameter integer VC0_TOTAL_CREDITS_CH = 31;
    parameter integer VC0_TOTAL_CREDITS_NPH = 12;
    parameter integer VC0_TOTAL_CREDITS_PD = 288;
    parameter integer VC0_TOTAL_CREDITS_PH = 32;
    parameter integer VC0_TX_LASTPACKET = 31;
    parameter [11:0] VC_BASE_PTR = 12'h10C;
    parameter [15:0] VC_CAP_ID = 16'h0002;
    parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
    parameter VC_CAP_ON = "FALSE";
    parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
    parameter [3:0] VC_CAP_VERSION = 4'h1;
    parameter [15:0] VENDOR_ID = 16'h10EE;
    parameter [11:0] VSEC_BASE_PTR = 12'h160;
    parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
    parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
    parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
    parameter [15:0] VSEC_CAP_ID = 16'h000B;
    parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
    parameter [11:0] VSEC_CAP_NEXTPTR = 12'h000;
    parameter VSEC_CAP_ON = "FALSE";
    parameter [3:0] VSEC_CAP_VERSION = 4'h1;
    output CFGAERECRCCHECKEN;
    output CFGAERECRCGENEN;
    output CFGCOMMANDBUSMASTERENABLE;
    output CFGCOMMANDINTERRUPTDISABLE;
    output CFGCOMMANDIOENABLE;
    output CFGCOMMANDMEMENABLE;
    output CFGCOMMANDSERREN;
    output CFGDEVCONTROL2CPLTIMEOUTDIS;
    output CFGDEVCONTROLAUXPOWEREN;
    output CFGDEVCONTROLCORRERRREPORTINGEN;
    output CFGDEVCONTROLENABLERO;
    output CFGDEVCONTROLEXTTAGEN;
    output CFGDEVCONTROLFATALERRREPORTINGEN;
    output CFGDEVCONTROLNONFATALREPORTINGEN;
    output CFGDEVCONTROLNOSNOOPEN;
    output CFGDEVCONTROLPHANTOMEN;
    output CFGDEVCONTROLURERRREPORTINGEN;
    output CFGDEVSTATUSCORRERRDETECTED;
    output CFGDEVSTATUSFATALERRDETECTED;
    output CFGDEVSTATUSNONFATALERRDETECTED;
    output CFGDEVSTATUSURDETECTED;
    output CFGERRAERHEADERLOGSETN;
    output CFGERRCPLRDYN;
    output CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFM;
    output CFGINTERRUPTRDYN;
    output CFGLINKCONTROLAUTOBANDWIDTHINTEN;
    output CFGLINKCONTROLBANDWIDTHINTEN;
    output CFGLINKCONTROLCLOCKPMEN;
    output CFGLINKCONTROLCOMMONCLOCK;
    output CFGLINKCONTROLEXTENDEDSYNC;
    output CFGLINKCONTROLHWAUTOWIDTHDIS;
    output CFGLINKCONTROLLINKDISABLE;
    output CFGLINKCONTROLRCB;
    output CFGLINKCONTROLRETRAINLINK;
    output CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
    output CFGLINKSTATUSBANDWITHSTATUS;
    output CFGLINKSTATUSDLLACTIVE;
    output CFGLINKSTATUSLINKTRAINING;
    output CFGMSGRECEIVED;
    output CFGMSGRECEIVEDASSERTINTA;
    output CFGMSGRECEIVEDASSERTINTB;
    output CFGMSGRECEIVEDASSERTINTC;
    output CFGMSGRECEIVEDASSERTINTD;
    output CFGMSGRECEIVEDDEASSERTINTA;
    output CFGMSGRECEIVEDDEASSERTINTB;
    output CFGMSGRECEIVEDDEASSERTINTC;
    output CFGMSGRECEIVEDDEASSERTINTD;
    output CFGMSGRECEIVEDERRCOR;
    output CFGMSGRECEIVEDERRFATAL;
    output CFGMSGRECEIVEDERRNONFATAL;
    output CFGMSGRECEIVEDPMASNAK;
    output CFGMSGRECEIVEDPMETO;
    output CFGMSGRECEIVEDPMETOACK;
    output CFGMSGRECEIVEDPMPME;
    output CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
    output CFGMSGRECEIVEDUNLOCK;
    output CFGPMCSRPMEEN;
    output CFGPMCSRPMESTATUS;
    output CFGPMRCVASREQL1N;
    output CFGPMRCVENTERL1N;
    output CFGPMRCVENTERL23N;
    output CFGPMRCVREQACKN;
    output CFGRDWRDONEN;
    output CFGSLOTCONTROLELECTROMECHILCTLPULSE;
    output CFGTRANSACTION;
    output CFGTRANSACTIONTYPE;
    output DBGSCLRA;
    output DBGSCLRB;
    output DBGSCLRC;
    output DBGSCLRD;
    output DBGSCLRE;
    output DBGSCLRF;
    output DBGSCLRG;
    output DBGSCLRH;
    output DBGSCLRI;
    output DBGSCLRJ;
    output DBGSCLRK;
    output DRPDRDY;
    output LL2BADDLLPERRN;
    output LL2BADTLPERRN;
    output LL2PROTOCOLERRN;
    output LL2REPLAYROERRN;
    output LL2REPLAYTOERRN;
    output LL2SUSPENDOKN;
    output LL2TFCINIT1SEQN;
    output LL2TFCINIT2SEQN;
    output LNKCLKEN;
    output MIMRXRCE;
    output MIMRXREN;
    output MIMRXWEN;
    output MIMTXRCE;
    output MIMTXREN;
    output MIMTXWEN;
    output PIPERX0POLARITY;
    output PIPERX1POLARITY;
    output PIPERX2POLARITY;
    output PIPERX3POLARITY;
    output PIPERX4POLARITY;
    output PIPERX5POLARITY;
    output PIPERX6POLARITY;
    output PIPERX7POLARITY;
    output PIPETX0COMPLIANCE;
    output PIPETX0ELECIDLE;
    output PIPETX1COMPLIANCE;
    output PIPETX1ELECIDLE;
    output PIPETX2COMPLIANCE;
    output PIPETX2ELECIDLE;
    output PIPETX3COMPLIANCE;
    output PIPETX3ELECIDLE;
    output PIPETX4COMPLIANCE;
    output PIPETX4ELECIDLE;
    output PIPETX5COMPLIANCE;
    output PIPETX5ELECIDLE;
    output PIPETX6COMPLIANCE;
    output PIPETX6ELECIDLE;
    output PIPETX7COMPLIANCE;
    output PIPETX7ELECIDLE;
    output PIPETXDEEMPH;
    output PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PL2LINKUPN;
    output PL2RECEIVERERRN;
    output PL2RECOVERYN;
    output PL2RXELECIDLE;
    output PL2SUSPENDOK;
    output PLLINKGEN2CAP;
    output PLLINKPARTNERGEN2SUPPORTED;
    output PLLINKUPCFGCAP;
    output PLPHYLNKUPN;
    output PLRECEIVEDHOTRST;
    output PLSELLNKRATE;
    output RECEIVEDFUNCLVLRSTN;
    output TL2ASPMSUSPENDCREDITCHECKOKN;
    output TL2ASPMSUSPENDREQN;
    output TL2PPMSUSPENDOKN;
    output TRNLNKUPN;
    output TRNRDLLPSRCRDYN;
    output TRNRECRCERRN;
    output TRNREOFN;
    output TRNRERRFWDN;
    output TRNRREMN;
    output TRNRSOFN;
    output TRNRSRCDSCN;
    output TRNRSRCRDYN;
    output TRNTCFGREQN;
    output TRNTDLLPDSTRDYN;
    output TRNTDSTRDYN;
    output TRNTERRDROPN;
    output USERRSTN;
    output [11:0] DBGVECC;
    output [11:0] PLDBGVEC;
    output [11:0] TRNFCCPLD;
    output [11:0] TRNFCNPD;
    output [11:0] TRNFCPD;
    output [12:0] MIMRXRADDR;
    output [12:0] MIMRXWADDR;
    output [12:0] MIMTXRADDR;
    output [12:0] MIMTXWADDR;
    output [15:0] CFGMSGDATA;
    output [15:0] DRPDO;
    output [15:0] PIPETX0DATA;
    output [15:0] PIPETX1DATA;
    output [15:0] PIPETX2DATA;
    output [15:0] PIPETX3DATA;
    output [15:0] PIPETX4DATA;
    output [15:0] PIPETX5DATA;
    output [15:0] PIPETX6DATA;
    output [15:0] PIPETX7DATA;
    output [1:0] CFGLINKCONTROLASPMCONTROL;
    output [1:0] CFGLINKSTATUSCURRENTSPEED;
    output [1:0] CFGPMCSRPOWERSTATE;
    output [1:0] PIPETX0CHARISK;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX1CHARISK;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX2CHARISK;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX3CHARISK;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX4CHARISK;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX5CHARISK;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX6CHARISK;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX7CHARISK;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PLLANEREVERSALMODE;
    output [1:0] PLRXPMSTATE;
    output [1:0] PLSELLNKWIDTH;
    output [2:0] CFGDEVCONTROLMAXPAYLOAD;
    output [2:0] CFGDEVCONTROLMAXREADREQ;
    output [2:0] CFGINTERRUPTMMENABLE;
    output [2:0] CFGPCIELINKSTATE;
    output [2:0] PIPETXMARGIN;
    output [2:0] PLINITIALLINKWIDTH;
    output [2:0] PLTXPMSTATE;
    output [31:0] CFGDO;
    output [31:0] TRNRDLLPDATA;
    output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL;
    output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH;
    output [5:0] PLLTSSMSTATE;
    output [5:0] TRNTBUFAV;
    output [63:0] DBGVECA;
    output [63:0] DBGVECB;
    output [63:0] TRNRD;
    output [67:0] MIMRXWDATA;
    output [68:0] MIMTXWDATA;
    output [6:0] CFGTRANSACTIONADDR;
    output [6:0] CFGVCTCVCMAP;
    output [6:0] TRNRBARHITN;
    output [7:0] CFGINTERRUPTDO;
    output [7:0] TRNFCCPLH;
    output [7:0] TRNFCNPH;
    output [7:0] TRNFCPH;
    input CFGERRACSN;
    input CFGERRCORN;
    input CFGERRCPLABORTN;
    input CFGERRCPLTIMEOUTN;
    input CFGERRCPLUNEXPECTN;
    input CFGERRECRCN;
    input CFGERRLOCKEDN;
    input CFGERRPOSTEDN;
    input CFGERRURN;
    input CFGINTERRUPTASSERTN;
    input CFGINTERRUPTN;
    input CFGPMDIRECTASPML1N;
    input CFGPMSENDPMACKN;
    input CFGPMSENDPMETON;
    input CFGPMSENDPMNAKN;
    input CFGPMTURNOFFOKN;
    input CFGPMWAKEN;
    input CFGRDENN;
    input CFGTRNPENDINGN;
    input CFGWRENN;
    input CFGWRREADONLYN;
    input CFGWRRW1CASRWN;
    input CMRSTN;
    input CMSTICKYRSTN;
    input DBGSUBMODE;
    input DLRSTN;
    input DRPCLK;
    input DRPDEN;
    input DRPDWE;
    input FUNCLVLRSTN;
    input LL2SENDASREQL1N;
    input LL2SENDENTERL1N;
    input LL2SENDENTERL23N;
    input LL2SUSPENDNOWN;
    input LL2TLPRCVN;
    input PIPECLK;
    input PIPERX0CHANISALIGNED;
    input PIPERX0ELECIDLE;
    input PIPERX0PHYSTATUS;
    input PIPERX0VALID;
    input PIPERX1CHANISALIGNED;
    input PIPERX1ELECIDLE;
    input PIPERX1PHYSTATUS;
    input PIPERX1VALID;
    input PIPERX2CHANISALIGNED;
    input PIPERX2ELECIDLE;
    input PIPERX2PHYSTATUS;
    input PIPERX2VALID;
    input PIPERX3CHANISALIGNED;
    input PIPERX3ELECIDLE;
    input PIPERX3PHYSTATUS;
    input PIPERX3VALID;
    input PIPERX4CHANISALIGNED;
    input PIPERX4ELECIDLE;
    input PIPERX4PHYSTATUS;
    input PIPERX4VALID;
    input PIPERX5CHANISALIGNED;
    input PIPERX5ELECIDLE;
    input PIPERX5PHYSTATUS;
    input PIPERX5VALID;
    input PIPERX6CHANISALIGNED;
    input PIPERX6ELECIDLE;
    input PIPERX6PHYSTATUS;
    input PIPERX6VALID;
    input PIPERX7CHANISALIGNED;
    input PIPERX7ELECIDLE;
    input PIPERX7PHYSTATUS;
    input PIPERX7VALID;
    input PLDIRECTEDLINKAUTON;
    input PLDIRECTEDLINKSPEED;
    input PLDOWNSTREAMDEEMPHSOURCE;
    input PLRSTN;
    input PLTRANSMITHOTRST;
    input PLUPSTREAMPREFERDEEMPH;
    input SYSRSTN;
    input TL2ASPMSUSPENDCREDITCHECKN;
    input TL2PPMSUSPENDREQN;
    input TLRSTN;
    input TRNRDSTRDYN;
    input TRNRNPOKN;
    input TRNTCFGGNTN;
    input TRNTDLLPSRCRDYN;
    input TRNTECRCGENN;
    input TRNTEOFN;
    input TRNTERRFWDN;
    input TRNTREMN;
    input TRNTSOFN;
    input TRNTSRCDSCN;
    input TRNTSRCRDYN;
    input TRNTSTRN;
    input USERCLK;
    input [127:0] CFGERRAERHEADERLOG;
    input [15:0] DRPDI;
    input [15:0] PIPERX0DATA;
    input [15:0] PIPERX1DATA;
    input [15:0] PIPERX2DATA;
    input [15:0] PIPERX3DATA;
    input [15:0] PIPERX4DATA;
    input [15:0] PIPERX5DATA;
    input [15:0] PIPERX6DATA;
    input [15:0] PIPERX7DATA;
    input [1:0] DBGMODE;
    input [1:0] PIPERX0CHARISK;
    input [1:0] PIPERX1CHARISK;
    input [1:0] PIPERX2CHARISK;
    input [1:0] PIPERX3CHARISK;
    input [1:0] PIPERX4CHARISK;
    input [1:0] PIPERX5CHARISK;
    input [1:0] PIPERX6CHARISK;
    input [1:0] PIPERX7CHARISK;
    input [1:0] PLDIRECTEDLINKCHANGE;
    input [1:0] PLDIRECTEDLINKWIDTH;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [2:0] PIPERX0STATUS;
    input [2:0] PIPERX1STATUS;
    input [2:0] PIPERX2STATUS;
    input [2:0] PIPERX3STATUS;
    input [2:0] PIPERX4STATUS;
    input [2:0] PIPERX5STATUS;
    input [2:0] PIPERX6STATUS;
    input [2:0] PIPERX7STATUS;
    input [2:0] PLDBGMODE;
    input [2:0] TRNFCSEL;
    input [31:0] CFGDI;
    input [31:0] TRNTDLLPDATA;
    input [3:0] CFGBYTEENN;
    input [47:0] CFGERRTLPCPLHEADER;
    input [4:0] CFGDSDEVICENUMBER;
    input [4:0] PL2DIRECTEDLSTATE;
    input [63:0] CFGDSN;
    input [63:0] TRNTD;
    input [67:0] MIMRXRDATA;
    input [68:0] MIMTXRDATA;
    input [7:0] CFGDSBUSNUMBER;
    input [7:0] CFGINTERRUPTDI;
    input [7:0] CFGPORTNUMBER;
    input [8:0] DRPDADDR;
    input [9:0] CFGDWADDR;
endmodule

module SYSMON (...);
    output BUSY;
    output DRDY;
    output EOC;
    output EOS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output OT;
    output [15:0] DO;
    output [2:0] ALM;
    output [4:0] CHANNEL;
    input CONVST;
    input CONVSTCLK;
    input DCLK;
    input DEN;
    input DWE;
    input RESET;
    input VN;
    input VP;
    input [15:0] DI;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input [6:0] DADDR;
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0800;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter SIM_DEVICE = "VIRTEX5";
    parameter SIM_MONITOR_FILE = "design.txt";
endmodule

module DSP48E1 (...);
    parameter integer ACASCREG = 1;
    parameter integer ADREG = 1;
    parameter integer ALUMODEREG = 1;
    parameter integer AREG = 1;
    parameter AUTORESET_PATDET = "NO_RESET";
    parameter A_INPUT = "DIRECT";
    parameter integer BCASCREG = 1;
    parameter integer BREG = 1;
    parameter B_INPUT = "DIRECT";
    parameter integer CARRYINREG = 1;
    parameter integer CARRYINSELREG = 1;
    parameter integer CREG = 1;
    parameter integer DREG = 1;
    parameter integer INMODEREG = 1;
    parameter integer MREG = 1;
    parameter integer OPMODEREG = 1;
    parameter integer PREG = 1;
    parameter SEL_MASK = "MASK";
    parameter SEL_PATTERN = "PATTERN";
    parameter USE_DPORT = "FALSE";
    parameter USE_MULT = "MULTIPLY";
    parameter USE_PATTERN_DETECT = "NO_PATDET";
    parameter USE_SIMD = "ONE48";
    parameter [47:0] MASK = 48'h3FFFFFFFFFFF;
    parameter [47:0] PATTERN = 48'h000000000000;
    parameter [3:0] IS_ALUMODE_INVERTED = 4'b0;
    parameter [0:0] IS_CARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [4:0] IS_INMODE_INVERTED = 5'b0;
    parameter [6:0] IS_OPMODE_INVERTED = 7'b0;
    output [29:0] ACOUT;
    output [17:0] BCOUT;
    output CARRYCASCOUT;
    output [3:0] CARRYOUT;
    output MULTSIGNOUT;
    output OVERFLOW;
    output [47:0] P;
    output PATTERNBDETECT;
    output PATTERNDETECT;
    output [47:0] PCOUT;
    output UNDERFLOW;
    input [29:0] A;
    input [29:0] ACIN;
    input [3:0] ALUMODE;
    input [17:0] B;
    input [17:0] BCIN;
    input [47:0] C;
    input CARRYCASCIN;
    input CARRYIN;
    input [2:0] CARRYINSEL;
    input CEA1;
    input CEA2;
    input CEAD;
    input CEALUMODE;
    input CEB1;
    input CEB2;
    input CEC;
    input CECARRYIN;
    input CECTRL;
    input CED;
    input CEINMODE;
    input CEM;
    input CEP;
    (* clkbuf_sink *)
    input CLK;
    input [24:0] D;
    input [4:0] INMODE;
    input MULTSIGNIN;
    input [6:0] OPMODE;
    input [47:0] PCIN;
    input RSTA;
    input RSTALLCARRYIN;
    input RSTALUMODE;
    input RSTB;
    input RSTC;
    input RSTCTRL;
    input RSTD;
    input RSTINMODE;
    input RSTM;
    input RSTP;
endmodule

module BUFGCE (...);
    parameter CE_TYPE = "SYNC";
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    input CE;
    input I;
endmodule

module BUFGCE_1 (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input I;
endmodule

module BUFGMUX (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_1 (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_CTRL (...);
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFH (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFIO (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFIODQS (...);
    parameter DQSMASK_ENABLE = "FALSE";
    (* clkbuf_driver *)
    output O;
    input DQSMASK;
    input I;
endmodule

module BUFR (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input CLR;
    input I;
    parameter BUFR_DIVIDE = "BYPASS";
    parameter SIM_DEVICE = "7SERIES";
endmodule

module IBUFDS_GTXE1 (...);
    parameter CLKCM_CFG = "TRUE";
    parameter CLKRCV_TRST = "TRUE";
    parameter [9:0] REFCLKOUT_DLY = 10'b0000000000;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module MMCM_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter CLOCK_HOLD = "FALSE";
    parameter COMPENSATION = "ZHOLD";
    parameter STARTUP_WAIT = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter real VCOCLK_FREQ_MAX = 1600.0;
    parameter real VCOCLK_FREQ_MIN = 600.0;
    parameter real CLKIN_FREQ_MAX = 800.0;
    parameter real CLKIN_FREQ_MIN = 10.0;
    parameter real CLKPFD_FREQ_MAX = 550.0;
    parameter real CLKPFD_FREQ_MIN = 10.0;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output DRDY;
    output LOCKED;
    output PSDONE;
    output [15:0] DO;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    input CLKINSEL;
    input DCLK;
    input DEN;
    input DWE;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input PWRDWN;
    input RST;
    input [15:0] DI;
    input [6:0] DADDR;
endmodule

module MMCM_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLOCK_HOLD = "FALSE";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

(* keep *)
module BSCAN_VIRTEX6 (...);
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
    parameter DISABLE_JTAG = "FALSE";
    parameter integer JTAG_CHAIN = 1;
endmodule

(* keep *)
module CAPTURE_VIRTEX6 (...);
    input CAP;
    input CLK;
    parameter ONESHOT = "TRUE";
endmodule

module DNA_PORT (...);
    parameter [56:0] SIM_DNA_VALUE = 57'h0;
    output DOUT;
    input CLK;
    input DIN;
    input READ;
    input SHIFT;
endmodule

module EFUSE_USR (...);
    parameter [31:0] SIM_EFUSE_VALUE = 32'h00000000;
    output [31:0] EFUSEUSR;
endmodule

module FRAME_ECC_VIRTEX6 (...);
    parameter FARSRC = "EFAR";
    parameter FRAME_RBT_IN_FILENAME = "NONE";
    output CRCERROR;
    output ECCERROR;
    output ECCERRORSINGLE;
    output SYNDROMEVALID;
    output [12:0] SYNDROME;
    output [23:0] FAR;
    output [4:0] SYNBIT;
    output [6:0] SYNWORD;
endmodule

(* keep *)
module ICAP_VIRTEX6 (...);
    parameter [31:0] DEVICE_ID = 32'h04244093;
    parameter ICAP_WIDTH = "X8";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output BUSY;
    output [31:0] O;
    input CLK;
    input CSB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module STARTUP_VIRTEX6 (...);
    parameter PROG_USR = "FALSE";
    output CFGCLK;
    output CFGMCLK;
    output DINSPI;
    output EOS;
    output PREQ;
    output TCKSPI;
    input CLK;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

module USR_ACCESS_VIRTEX6 (...);
    output CFGCLK;
    output [31:0] DATA;
    output DATAVALID;
endmodule

(* keep *)
module DCIRESET (...);
    output LOCKED;
    input RST;
endmodule

module GTHE1_QUAD (...);
    parameter [15:0] BER_CONST_PTRN0 = 16'h0000;
    parameter [15:0] BER_CONST_PTRN1 = 16'h0000;
    parameter [15:0] BUFFER_CONFIG_LANE0 = 16'h4004;
    parameter [15:0] BUFFER_CONFIG_LANE1 = 16'h4004;
    parameter [15:0] BUFFER_CONFIG_LANE2 = 16'h4004;
    parameter [15:0] BUFFER_CONFIG_LANE3 = 16'h4004;
    parameter [15:0] DFE_TRAIN_CTRL_LANE0 = 16'h0000;
    parameter [15:0] DFE_TRAIN_CTRL_LANE1 = 16'h0000;
    parameter [15:0] DFE_TRAIN_CTRL_LANE2 = 16'h0000;
    parameter [15:0] DFE_TRAIN_CTRL_LANE3 = 16'h0000;
    parameter [15:0] DLL_CFG0 = 16'h8202;
    parameter [15:0] DLL_CFG1 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEKR_LD_COEFF_UPD_LANE3 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEKR_LP_COEFF_UPD_LANE3 = 16'h0000;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE0 = 16'h0002;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE1 = 16'h0002;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE2 = 16'h0002;
    parameter [15:0] E10GBASEKR_PMA_CTRL_LANE3 = 16'h0002;
    parameter [15:0] E10GBASEKX_CTRL_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEKX_CTRL_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEKX_CTRL_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEKX_CTRL_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_CFG_LANE0 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_CFG_LANE1 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_CFG_LANE2 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_CFG_LANE3 = 16'h070C;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE0 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE1 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE2 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA0_LANE3 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA1_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA2_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDA3_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE0 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE1 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE2 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB0_LANE3 = 16'h0001;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB1_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB2_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_SEEDB3_LANE3 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE0 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE1 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE2 = 16'h0000;
    parameter [15:0] E10GBASER_PCS_TEST_CTRL_LANE3 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE0 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE1 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE2 = 16'h0000;
    parameter [15:0] E10GBASEX_PCS_TSTCTRL_LANE3 = 16'h0000;
    parameter [15:0] GLBL0_NOISE_CTRL = 16'hF0B8;
    parameter [15:0] GLBL_AMON_SEL = 16'h0000;
    parameter [15:0] GLBL_DMON_SEL = 16'h0200;
    parameter [15:0] GLBL_PWR_CTRL = 16'h0000;
    parameter [0:0] GTH_CFG_PWRUP_LANE0 = 1'b1;
    parameter [0:0] GTH_CFG_PWRUP_LANE1 = 1'b1;
    parameter [0:0] GTH_CFG_PWRUP_LANE2 = 1'b1;
    parameter [0:0] GTH_CFG_PWRUP_LANE3 = 1'b1;
    parameter [15:0] LANE_AMON_SEL = 16'h00F0;
    parameter [15:0] LANE_DMON_SEL = 16'h0000;
    parameter [15:0] LANE_LNK_CFGOVRD = 16'h0000;
    parameter [15:0] LANE_PWR_CTRL_LANE0 = 16'h0400;
    parameter [15:0] LANE_PWR_CTRL_LANE1 = 16'h0400;
    parameter [15:0] LANE_PWR_CTRL_LANE2 = 16'h0400;
    parameter [15:0] LANE_PWR_CTRL_LANE3 = 16'h0400;
    parameter [15:0] LNK_TRN_CFG_LANE0 = 16'h0000;
    parameter [15:0] LNK_TRN_CFG_LANE1 = 16'h0000;
    parameter [15:0] LNK_TRN_CFG_LANE2 = 16'h0000;
    parameter [15:0] LNK_TRN_CFG_LANE3 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE0 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE1 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE2 = 16'h0000;
    parameter [15:0] LNK_TRN_COEFF_REQ_LANE3 = 16'h0000;
    parameter [15:0] MISC_CFG = 16'h0008;
    parameter [15:0] MODE_CFG1 = 16'h0000;
    parameter [15:0] MODE_CFG2 = 16'h0000;
    parameter [15:0] MODE_CFG3 = 16'h0000;
    parameter [15:0] MODE_CFG4 = 16'h0000;
    parameter [15:0] MODE_CFG5 = 16'h0000;
    parameter [15:0] MODE_CFG6 = 16'h0000;
    parameter [15:0] MODE_CFG7 = 16'h0000;
    parameter [15:0] PCS_ABILITY_LANE0 = 16'h0010;
    parameter [15:0] PCS_ABILITY_LANE1 = 16'h0010;
    parameter [15:0] PCS_ABILITY_LANE2 = 16'h0010;
    parameter [15:0] PCS_ABILITY_LANE3 = 16'h0010;
    parameter [15:0] PCS_CTRL1_LANE0 = 16'h2040;
    parameter [15:0] PCS_CTRL1_LANE1 = 16'h2040;
    parameter [15:0] PCS_CTRL1_LANE2 = 16'h2040;
    parameter [15:0] PCS_CTRL1_LANE3 = 16'h2040;
    parameter [15:0] PCS_CTRL2_LANE0 = 16'h0000;
    parameter [15:0] PCS_CTRL2_LANE1 = 16'h0000;
    parameter [15:0] PCS_CTRL2_LANE2 = 16'h0000;
    parameter [15:0] PCS_CTRL2_LANE3 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_0_LANE0 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_0_LANE1 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_0_LANE2 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_0_LANE3 = 16'h1116;
    parameter [15:0] PCS_MISC_CFG_1_LANE0 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_1_LANE1 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_1_LANE2 = 16'h0000;
    parameter [15:0] PCS_MISC_CFG_1_LANE3 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE0 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE1 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE2 = 16'h0000;
    parameter [15:0] PCS_MODE_LANE3 = 16'h0000;
    parameter [15:0] PCS_RESET_1_LANE0 = 16'h0002;
    parameter [15:0] PCS_RESET_1_LANE1 = 16'h0002;
    parameter [15:0] PCS_RESET_1_LANE2 = 16'h0002;
    parameter [15:0] PCS_RESET_1_LANE3 = 16'h0002;
    parameter [15:0] PCS_RESET_LANE0 = 16'h0000;
    parameter [15:0] PCS_RESET_LANE1 = 16'h0000;
    parameter [15:0] PCS_RESET_LANE2 = 16'h0000;
    parameter [15:0] PCS_RESET_LANE3 = 16'h0000;
    parameter [15:0] PCS_TYPE_LANE0 = 16'h002C;
    parameter [15:0] PCS_TYPE_LANE1 = 16'h002C;
    parameter [15:0] PCS_TYPE_LANE2 = 16'h002C;
    parameter [15:0] PCS_TYPE_LANE3 = 16'h002C;
    parameter [15:0] PLL_CFG0 = 16'h95DF;
    parameter [15:0] PLL_CFG1 = 16'h81C0;
    parameter [15:0] PLL_CFG2 = 16'h0424;
    parameter [15:0] PMA_CTRL1_LANE0 = 16'h0000;
    parameter [15:0] PMA_CTRL1_LANE1 = 16'h0000;
    parameter [15:0] PMA_CTRL1_LANE2 = 16'h0000;
    parameter [15:0] PMA_CTRL1_LANE3 = 16'h0000;
    parameter [15:0] PMA_CTRL2_LANE0 = 16'h000B;
    parameter [15:0] PMA_CTRL2_LANE1 = 16'h000B;
    parameter [15:0] PMA_CTRL2_LANE2 = 16'h000B;
    parameter [15:0] PMA_CTRL2_LANE3 = 16'h000B;
    parameter [15:0] PMA_LPBK_CTRL_LANE0 = 16'h0004;
    parameter [15:0] PMA_LPBK_CTRL_LANE1 = 16'h0004;
    parameter [15:0] PMA_LPBK_CTRL_LANE2 = 16'h0004;
    parameter [15:0] PMA_LPBK_CTRL_LANE3 = 16'h0004;
    parameter [15:0] PRBS_BER_CFG0_LANE0 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG0_LANE1 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG0_LANE2 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG0_LANE3 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE0 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE1 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE2 = 16'h0000;
    parameter [15:0] PRBS_BER_CFG1_LANE3 = 16'h0000;
    parameter [15:0] PRBS_CFG_LANE0 = 16'h000A;
    parameter [15:0] PRBS_CFG_LANE1 = 16'h000A;
    parameter [15:0] PRBS_CFG_LANE2 = 16'h000A;
    parameter [15:0] PRBS_CFG_LANE3 = 16'h000A;
    parameter [15:0] PTRN_CFG0_LSB = 16'h5555;
    parameter [15:0] PTRN_CFG0_MSB = 16'h5555;
    parameter [15:0] PTRN_LEN_CFG = 16'h001F;
    parameter [15:0] PWRUP_DLY = 16'h0000;
    parameter [15:0] RX_AEQ_VAL0_LANE0 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL0_LANE1 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL0_LANE2 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL0_LANE3 = 16'h03C0;
    parameter [15:0] RX_AEQ_VAL1_LANE0 = 16'h0000;
    parameter [15:0] RX_AEQ_VAL1_LANE1 = 16'h0000;
    parameter [15:0] RX_AEQ_VAL1_LANE2 = 16'h0000;
    parameter [15:0] RX_AEQ_VAL1_LANE3 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE0 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE1 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE2 = 16'h0000;
    parameter [15:0] RX_AGC_CTRL_LANE3 = 16'h0000;
    parameter [15:0] RX_CDR_CTRL0_LANE0 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL0_LANE1 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL0_LANE2 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL0_LANE3 = 16'h0005;
    parameter [15:0] RX_CDR_CTRL1_LANE0 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL1_LANE1 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL1_LANE2 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL1_LANE3 = 16'h4200;
    parameter [15:0] RX_CDR_CTRL2_LANE0 = 16'h2000;
    parameter [15:0] RX_CDR_CTRL2_LANE1 = 16'h2000;
    parameter [15:0] RX_CDR_CTRL2_LANE2 = 16'h2000;
    parameter [15:0] RX_CDR_CTRL2_LANE3 = 16'h2000;
    parameter [15:0] RX_CFG0_LANE0 = 16'h0500;
    parameter [15:0] RX_CFG0_LANE1 = 16'h0500;
    parameter [15:0] RX_CFG0_LANE2 = 16'h0500;
    parameter [15:0] RX_CFG0_LANE3 = 16'h0500;
    parameter [15:0] RX_CFG1_LANE0 = 16'h821F;
    parameter [15:0] RX_CFG1_LANE1 = 16'h821F;
    parameter [15:0] RX_CFG1_LANE2 = 16'h821F;
    parameter [15:0] RX_CFG1_LANE3 = 16'h821F;
    parameter [15:0] RX_CFG2_LANE0 = 16'h1001;
    parameter [15:0] RX_CFG2_LANE1 = 16'h1001;
    parameter [15:0] RX_CFG2_LANE2 = 16'h1001;
    parameter [15:0] RX_CFG2_LANE3 = 16'h1001;
    parameter [15:0] RX_CTLE_CTRL_LANE0 = 16'h008F;
    parameter [15:0] RX_CTLE_CTRL_LANE1 = 16'h008F;
    parameter [15:0] RX_CTLE_CTRL_LANE2 = 16'h008F;
    parameter [15:0] RX_CTLE_CTRL_LANE3 = 16'h008F;
    parameter [15:0] RX_CTRL_OVRD_LANE0 = 16'h000C;
    parameter [15:0] RX_CTRL_OVRD_LANE1 = 16'h000C;
    parameter [15:0] RX_CTRL_OVRD_LANE2 = 16'h000C;
    parameter [15:0] RX_CTRL_OVRD_LANE3 = 16'h000C;
    parameter integer RX_FABRIC_WIDTH0 = 6466;
    parameter integer RX_FABRIC_WIDTH1 = 6466;
    parameter integer RX_FABRIC_WIDTH2 = 6466;
    parameter integer RX_FABRIC_WIDTH3 = 6466;
    parameter [15:0] RX_LOOP_CTRL_LANE0 = 16'h007F;
    parameter [15:0] RX_LOOP_CTRL_LANE1 = 16'h007F;
    parameter [15:0] RX_LOOP_CTRL_LANE2 = 16'h007F;
    parameter [15:0] RX_LOOP_CTRL_LANE3 = 16'h007F;
    parameter [15:0] RX_MVAL0_LANE0 = 16'h0000;
    parameter [15:0] RX_MVAL0_LANE1 = 16'h0000;
    parameter [15:0] RX_MVAL0_LANE2 = 16'h0000;
    parameter [15:0] RX_MVAL0_LANE3 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE0 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE1 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE2 = 16'h0000;
    parameter [15:0] RX_MVAL1_LANE3 = 16'h0000;
    parameter [15:0] RX_P0S_CTRL = 16'h1206;
    parameter [15:0] RX_P0_CTRL = 16'h11F0;
    parameter [15:0] RX_P1_CTRL = 16'h120F;
    parameter [15:0] RX_P2_CTRL = 16'h0E0F;
    parameter [15:0] RX_PI_CTRL0 = 16'hD2F0;
    parameter [15:0] RX_PI_CTRL1 = 16'h0080;
    parameter integer SIM_GTHRESET_SPEEDUP = 1;
    parameter SIM_VERSION = "1.0";
    parameter [15:0] SLICE_CFG = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_0_LANE01 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_0_LANE23 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_1_LANE01 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_1_LANE23 = 16'h0000;
    parameter [15:0] SLICE_NOISE_CTRL_2_LANE01 = 16'h7FFF;
    parameter [15:0] SLICE_NOISE_CTRL_2_LANE23 = 16'h7FFF;
    parameter [15:0] SLICE_TX_RESET_LANE01 = 16'h0000;
    parameter [15:0] SLICE_TX_RESET_LANE23 = 16'h0000;
    parameter [15:0] TERM_CTRL_LANE0 = 16'h5007;
    parameter [15:0] TERM_CTRL_LANE1 = 16'h5007;
    parameter [15:0] TERM_CTRL_LANE2 = 16'h5007;
    parameter [15:0] TERM_CTRL_LANE3 = 16'h5007;
    parameter [15:0] TX_CFG0_LANE0 = 16'h203D;
    parameter [15:0] TX_CFG0_LANE1 = 16'h203D;
    parameter [15:0] TX_CFG0_LANE2 = 16'h203D;
    parameter [15:0] TX_CFG0_LANE3 = 16'h203D;
    parameter [15:0] TX_CFG1_LANE0 = 16'h0F00;
    parameter [15:0] TX_CFG1_LANE1 = 16'h0F00;
    parameter [15:0] TX_CFG1_LANE2 = 16'h0F00;
    parameter [15:0] TX_CFG1_LANE3 = 16'h0F00;
    parameter [15:0] TX_CFG2_LANE0 = 16'h0081;
    parameter [15:0] TX_CFG2_LANE1 = 16'h0081;
    parameter [15:0] TX_CFG2_LANE2 = 16'h0081;
    parameter [15:0] TX_CFG2_LANE3 = 16'h0081;
    parameter [15:0] TX_CLK_SEL0_LANE0 = 16'h2121;
    parameter [15:0] TX_CLK_SEL0_LANE1 = 16'h2121;
    parameter [15:0] TX_CLK_SEL0_LANE2 = 16'h2121;
    parameter [15:0] TX_CLK_SEL0_LANE3 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE0 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE1 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE2 = 16'h2121;
    parameter [15:0] TX_CLK_SEL1_LANE3 = 16'h2121;
    parameter [15:0] TX_DISABLE_LANE0 = 16'h0000;
    parameter [15:0] TX_DISABLE_LANE1 = 16'h0000;
    parameter [15:0] TX_DISABLE_LANE2 = 16'h0000;
    parameter [15:0] TX_DISABLE_LANE3 = 16'h0000;
    parameter integer TX_FABRIC_WIDTH0 = 6466;
    parameter integer TX_FABRIC_WIDTH1 = 6466;
    parameter integer TX_FABRIC_WIDTH2 = 6466;
    parameter integer TX_FABRIC_WIDTH3 = 6466;
    parameter [15:0] TX_P0P0S_CTRL = 16'h060C;
    parameter [15:0] TX_P1P2_CTRL = 16'h0C39;
    parameter [15:0] TX_PREEMPH_LANE0 = 16'h00A1;
    parameter [15:0] TX_PREEMPH_LANE1 = 16'h00A1;
    parameter [15:0] TX_PREEMPH_LANE2 = 16'h00A1;
    parameter [15:0] TX_PREEMPH_LANE3 = 16'h00A1;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE0 = 16'h0060;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE1 = 16'h0060;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE2 = 16'h0060;
    parameter [15:0] TX_PWR_RATE_OVRD_LANE3 = 16'h0060;
    output DRDY;
    output GTHINITDONE;
    output MGMTPCSRDACK;
    output RXCTRLACK0;
    output RXCTRLACK1;
    output RXCTRLACK2;
    output RXCTRLACK3;
    output RXDATATAP0;
    output RXDATATAP1;
    output RXDATATAP2;
    output RXDATATAP3;
    output RXPCSCLKSMPL0;
    output RXPCSCLKSMPL1;
    output RXPCSCLKSMPL2;
    output RXPCSCLKSMPL3;
    output RXUSERCLKOUT0;
    output RXUSERCLKOUT1;
    output RXUSERCLKOUT2;
    output RXUSERCLKOUT3;
    output TSTPATH;
    output TSTREFCLKFAB;
    output TSTREFCLKOUT;
    output TXCTRLACK0;
    output TXCTRLACK1;
    output TXCTRLACK2;
    output TXCTRLACK3;
    output TXDATATAP10;
    output TXDATATAP11;
    output TXDATATAP12;
    output TXDATATAP13;
    output TXDATATAP20;
    output TXDATATAP21;
    output TXDATATAP22;
    output TXDATATAP23;
    output TXN0;
    output TXN1;
    output TXN2;
    output TXN3;
    output TXP0;
    output TXP1;
    output TXP2;
    output TXP3;
    output TXPCSCLKSMPL0;
    output TXPCSCLKSMPL1;
    output TXPCSCLKSMPL2;
    output TXPCSCLKSMPL3;
    output TXUSERCLKOUT0;
    output TXUSERCLKOUT1;
    output TXUSERCLKOUT2;
    output TXUSERCLKOUT3;
    output [15:0] DRPDO;
    output [15:0] MGMTPCSRDDATA;
    output [63:0] RXDATA0;
    output [63:0] RXDATA1;
    output [63:0] RXDATA2;
    output [63:0] RXDATA3;
    output [7:0] RXCODEERR0;
    output [7:0] RXCODEERR1;
    output [7:0] RXCODEERR2;
    output [7:0] RXCODEERR3;
    output [7:0] RXCTRL0;
    output [7:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [7:0] RXDISPERR0;
    output [7:0] RXDISPERR1;
    output [7:0] RXDISPERR2;
    output [7:0] RXDISPERR3;
    output [7:0] RXVALID0;
    output [7:0] RXVALID1;
    output [7:0] RXVALID2;
    output [7:0] RXVALID3;
    input DCLK;
    input DEN;
    input DFETRAINCTRL0;
    input DFETRAINCTRL1;
    input DFETRAINCTRL2;
    input DFETRAINCTRL3;
    input DISABLEDRP;
    input DWE;
    input GTHINIT;
    input GTHRESET;
    input GTHX2LANE01;
    input GTHX2LANE23;
    input GTHX4LANE;
    input MGMTPCSREGRD;
    input MGMTPCSREGWR;
    input POWERDOWN0;
    input POWERDOWN1;
    input POWERDOWN2;
    input POWERDOWN3;
    input REFCLK;
    input RXBUFRESET0;
    input RXBUFRESET1;
    input RXBUFRESET2;
    input RXBUFRESET3;
    input RXENCOMMADET0;
    input RXENCOMMADET1;
    input RXENCOMMADET2;
    input RXENCOMMADET3;
    input RXN0;
    input RXN1;
    input RXN2;
    input RXN3;
    input RXP0;
    input RXP1;
    input RXP2;
    input RXP3;
    input RXPOLARITY0;
    input RXPOLARITY1;
    input RXPOLARITY2;
    input RXPOLARITY3;
    input RXSLIP0;
    input RXSLIP1;
    input RXSLIP2;
    input RXSLIP3;
    input RXUSERCLKIN0;
    input RXUSERCLKIN1;
    input RXUSERCLKIN2;
    input RXUSERCLKIN3;
    input TXBUFRESET0;
    input TXBUFRESET1;
    input TXBUFRESET2;
    input TXBUFRESET3;
    input TXDEEMPH0;
    input TXDEEMPH1;
    input TXDEEMPH2;
    input TXDEEMPH3;
    input TXUSERCLKIN0;
    input TXUSERCLKIN1;
    input TXUSERCLKIN2;
    input TXUSERCLKIN3;
    input [15:0] DADDR;
    input [15:0] DI;
    input [15:0] MGMTPCSREGADDR;
    input [15:0] MGMTPCSWRDATA;
    input [1:0] RXPOWERDOWN0;
    input [1:0] RXPOWERDOWN1;
    input [1:0] RXPOWERDOWN2;
    input [1:0] RXPOWERDOWN3;
    input [1:0] RXRATE0;
    input [1:0] RXRATE1;
    input [1:0] RXRATE2;
    input [1:0] RXRATE3;
    input [1:0] TXPOWERDOWN0;
    input [1:0] TXPOWERDOWN1;
    input [1:0] TXPOWERDOWN2;
    input [1:0] TXPOWERDOWN3;
    input [1:0] TXRATE0;
    input [1:0] TXRATE1;
    input [1:0] TXRATE2;
    input [1:0] TXRATE3;
    input [2:0] PLLREFCLKSEL;
    input [2:0] SAMPLERATE0;
    input [2:0] SAMPLERATE1;
    input [2:0] SAMPLERATE2;
    input [2:0] SAMPLERATE3;
    input [2:0] TXMARGIN0;
    input [2:0] TXMARGIN1;
    input [2:0] TXMARGIN2;
    input [2:0] TXMARGIN3;
    input [3:0] MGMTPCSLANESEL;
    input [4:0] MGMTPCSMMDADDR;
    input [5:0] PLLPCSCLKDIV;
    input [63:0] TXDATA0;
    input [63:0] TXDATA1;
    input [63:0] TXDATA2;
    input [63:0] TXDATA3;
    input [7:0] TXCTRL0;
    input [7:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [7:0] TXCTRL3;
    input [7:0] TXDATAMSB0;
    input [7:0] TXDATAMSB1;
    input [7:0] TXDATAMSB2;
    input [7:0] TXDATAMSB3;
endmodule

module GTXE1 (...);
    parameter AC_CAP_DIS = "TRUE";
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter [1:0] BGTEST_CFG = 2'b00;
    parameter [16:0] BIAS_CFG = 17'h00000;
    parameter [4:0] CDR_PH_ADJ_TIME = 5'b10100;
    parameter integer CHAN_BOND_1_MAX_SKEW = 7;
    parameter integer CHAN_BOND_2_MAX_SKEW = 1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0110111100;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100111100;
    parameter [4:0] CHAN_BOND_SEQ_2_CFG = 5'b00000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter integer CLK_COR_ADJ_LEN = 1;
    parameter integer CLK_COR_DET_LEN = 1;
    parameter CLK_COR_INSERT_IDLE_FLAG = "FALSE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter [1:0] CM_TRIM = 2'b01;
    parameter [9:0] COMMA_10B_ENABLE = 10'b1111111111;
    parameter COMMA_DOUBLE = "FALSE";
    parameter [3:0] COM_BURST_VAL = 4'b1111;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [4:0] DFE_CAL_TIME = 5'b01100;
    parameter [7:0] DFE_CFG = 8'b00011011;
    parameter [2:0] GEARBOX_ENDEC = 3'b000;
    parameter GEN_RXUSRCLK = "TRUE";
    parameter GEN_TXUSRCLK = "TRUE";
    parameter GTX_CFG_PWRUP = "TRUE";
    parameter [9:0] MCOMMA_10B_VALUE = 10'b1010000011;
    parameter MCOMMA_DETECT = "TRUE";
    parameter [2:0] OOBDETECT_THRESHOLD = 3'b011;
    parameter PCI_EXPRESS_MODE = "FALSE";
    parameter [9:0] PCOMMA_10B_VALUE = 10'b0101111100;
    parameter PCOMMA_DETECT = "TRUE";
    parameter PMA_CAS_CLK_EN = "FALSE";
    parameter [26:0] PMA_CDR_SCAN = 27'h640404C;
    parameter [75:0] PMA_CFG = 76'h0040000040000000003;
    parameter [6:0] PMA_RXSYNC_CFG = 7'h00;
    parameter [24:0] PMA_RX_CFG = 25'h05CE048;
    parameter [19:0] PMA_TX_CFG = 20'h00082;
    parameter [9:0] POWER_SAVE = 10'b0000110100;
    parameter RCV_TERM_GND = "FALSE";
    parameter RCV_TERM_VTTRX = "TRUE";
    parameter RXGEARBOX_USE = "FALSE";
    parameter [23:0] RXPLL_COM_CFG = 24'h21680A;
    parameter [7:0] RXPLL_CP_CFG = 8'h00;
    parameter integer RXPLL_DIVSEL45_FB = 5;
    parameter integer RXPLL_DIVSEL_FB = 2;
    parameter integer RXPLL_DIVSEL_OUT = 1;
    parameter integer RXPLL_DIVSEL_REF = 1;
    parameter [2:0] RXPLL_LKDET_CFG = 3'b111;
    parameter [0:0] RXPRBSERR_LOOPBACK = 1'b0;
    parameter RXRECCLK_CTRL = "RXRECCLKPCS";
    parameter [9:0] RXRECCLK_DLY = 10'b0000000000;
    parameter [15:0] RXUSRCLK_DLY = 16'h0000;
    parameter RX_BUFFER_USE = "TRUE";
    parameter integer RX_CLK25_DIVIDER = 6;
    parameter integer RX_DATA_WIDTH = 20;
    parameter RX_DECODE_SEQ_MATCH = "TRUE";
    parameter [3:0] RX_DLYALIGN_CTRINC = 4'b0100;
    parameter [4:0] RX_DLYALIGN_EDGESET = 5'b00110;
    parameter [3:0] RX_DLYALIGN_LPFINC = 4'b0111;
    parameter [2:0] RX_DLYALIGN_MONSEL = 3'b000;
    parameter [7:0] RX_DLYALIGN_OVRDSETTING = 8'b00000000;
    parameter RX_EN_IDLE_HOLD_CDR = "FALSE";
    parameter RX_EN_IDLE_HOLD_DFE = "TRUE";
    parameter RX_EN_IDLE_RESET_BUF = "TRUE";
    parameter RX_EN_IDLE_RESET_FR = "TRUE";
    parameter RX_EN_IDLE_RESET_PH = "TRUE";
    parameter RX_EN_MODE_RESET_BUF = "TRUE";
    parameter RX_EN_RATE_RESET_BUF = "TRUE";
    parameter RX_EN_REALIGN_RESET_BUF = "FALSE";
    parameter RX_EN_REALIGN_RESET_BUF2 = "FALSE";
    parameter [7:0] RX_EYE_OFFSET = 8'h4C;
    parameter [1:0] RX_EYE_SCANMODE = 2'b00;
    parameter RX_FIFO_ADDR_MODE = "FULL";
    parameter [3:0] RX_IDLE_HI_CNT = 4'b1000;
    parameter [3:0] RX_IDLE_LO_CNT = 4'b0000;
    parameter RX_LOSS_OF_SYNC_FSM = "FALSE";
    parameter integer RX_LOS_INVALID_INCR = 1;
    parameter integer RX_LOS_THRESHOLD = 4;
    parameter RX_OVERSAMPLE_MODE = "FALSE";
    parameter integer RX_SLIDE_AUTO_WAIT = 5;
    parameter RX_SLIDE_MODE = "OFF";
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COMSAS = 52;
    parameter integer SAS_MIN_COMSAS = 40;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter [2:0] SATA_IDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 7;
    parameter integer SATA_MAX_INIT = 22;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter integer SIM_GTXRESET_SPEEDUP = 1;
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter [2:0] SIM_RXREFCLK_SOURCE = 3'b000;
    parameter [2:0] SIM_TXREFCLK_SOURCE = 3'b000;
    parameter SIM_TX_ELEC_IDLE_LEVEL = "X";
    parameter SIM_VERSION = "2.0";
    parameter [4:0] TERMINATION_CTRL = 5'b10100;
    parameter TERMINATION_OVRD = "FALSE";
    parameter [11:0] TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] TRANS_TIME_NON_P2 = 8'h19;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [9:0] TRANS_TIME_TO_P2 = 10'h064;
    parameter [31:0] TST_ATTR = 32'h00000000;
    parameter TXDRIVE_LOOPBACK_HIZ = "FALSE";
    parameter TXDRIVE_LOOPBACK_PD = "FALSE";
    parameter TXGEARBOX_USE = "FALSE";
    parameter TXOUTCLK_CTRL = "TXOUTCLKPCS";
    parameter [9:0] TXOUTCLK_DLY = 10'b0000000000;
    parameter [23:0] TXPLL_COM_CFG = 24'h21680A;
    parameter [7:0] TXPLL_CP_CFG = 8'h00;
    parameter integer TXPLL_DIVSEL45_FB = 5;
    parameter integer TXPLL_DIVSEL_FB = 2;
    parameter integer TXPLL_DIVSEL_OUT = 1;
    parameter integer TXPLL_DIVSEL_REF = 1;
    parameter [2:0] TXPLL_LKDET_CFG = 3'b111;
    parameter [1:0] TXPLL_SATA = 2'b00;
    parameter TX_BUFFER_USE = "TRUE";
    parameter [5:0] TX_BYTECLK_CFG = 6'h00;
    parameter integer TX_CLK25_DIVIDER = 6;
    parameter TX_CLK_SOURCE = "RXPLL";
    parameter integer TX_DATA_WIDTH = 20;
    parameter [4:0] TX_DEEMPH_0 = 5'b11010;
    parameter [4:0] TX_DEEMPH_1 = 5'b10000;
    parameter [13:0] TX_DETECT_RX_CFG = 14'h1832;
    parameter [3:0] TX_DLYALIGN_CTRINC = 4'b0100;
    parameter [3:0] TX_DLYALIGN_LPFINC = 4'b0110;
    parameter [2:0] TX_DLYALIGN_MONSEL = 3'b000;
    parameter [7:0] TX_DLYALIGN_OVRDSETTING = 8'b10000000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter TX_EN_RATE_RESET_BUF = "TRUE";
    parameter [2:0] TX_IDLE_ASSERT_DELAY = 3'b100;
    parameter [2:0] TX_IDLE_DEASSERT_DELAY = 3'b010;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter TX_OVERSAMPLE_MODE = "FALSE";
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [1:0] TX_TDCC_CFG = 2'b11;
    parameter [5:0] TX_USRCLK_CFG = 6'h00;
    parameter TX_XCLK_SEL = "TXUSR";
    output COMFINISH;
    output COMINITDET;
    output COMSASDET;
    output COMWAKEDET;
    output DRDY;
    output PHYSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMMADET;
    output RXDATAVALID;
    output RXELECIDLE;
    output RXHEADERVALID;
    output RXOVERSAMPLEERR;
    output RXPLLLKDET;
    output RXPRBSERR;
    output RXRATEDONE;
    output RXRECCLK;
    output RXRECCLKPCS;
    output RXRESETDONE;
    output RXSTARTOFSEQ;
    output RXVALID;
    output TXGEARBOXREADY;
    output TXN;
    output TXOUTCLK;
    output TXOUTCLKPCS;
    output TXP;
    output TXPLLLKDET;
    output TXRATEDONE;
    output TXRESETDONE;
    output [15:0] DRPDO;
    output [1:0] MGTREFCLKFAB;
    output [1:0] RXLOSSOFSYNC;
    output [1:0] TXBUFSTATUS;
    output [2:0] DFESENSCAL;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXCLKCORCNT;
    output [2:0] RXHEADER;
    output [2:0] RXSTATUS;
    output [31:0] RXDATA;
    output [3:0] DFETAP3MONITOR;
    output [3:0] DFETAP4MONITOR;
    output [3:0] RXCHARISCOMMA;
    output [3:0] RXCHARISK;
    output [3:0] RXCHBONDO;
    output [3:0] RXDISPERR;
    output [3:0] RXNOTINTABLE;
    output [3:0] RXRUNDISP;
    output [3:0] TXKERR;
    output [3:0] TXRUNDISP;
    output [4:0] DFEEYEDACMON;
    output [4:0] DFETAP1MONITOR;
    output [4:0] DFETAP2MONITOR;
    output [5:0] DFECLKDLYADJMON;
    output [7:0] RXDLYALIGNMONITOR;
    output [7:0] TXDLYALIGNMONITOR;
    output [9:0] TSTOUT;
    input DCLK;
    input DEN;
    input DFEDLYOVRD;
    input DFETAPOVRD;
    input DWE;
    input GATERXELECIDLE;
    input GREFCLKRX;
    input GREFCLKTX;
    input GTXRXRESET;
    input GTXTXRESET;
    input IGNORESIGDET;
    input PERFCLKRX;
    input PERFCLKTX;
    input PLLRXRESET;
    input PLLTXRESET;
    input PRBSCNTRESET;
    input RXBUFRESET;
    input RXCDRRESET;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETUSE;
    input RXDEC8B10BUSE;
    input RXDLYALIGNDISABLE;
    input RXDLYALIGNMONENB;
    input RXDLYALIGNOVERRIDE;
    input RXDLYALIGNRESET;
    input RXDLYALIGNSWPPRECURB;
    input RXDLYALIGNUPDSW;
    input RXENCHANSYNC;
    input RXENMCOMMAALIGN;
    input RXENPCOMMAALIGN;
    input RXENPMAPHASEALIGN;
    input RXENSAMPLEALIGN;
    input RXGEARBOXSLIP;
    input RXN;
    input RXP;
    input RXPLLLKDETEN;
    input RXPLLPOWERDOWN;
    input RXPMASETPHASE;
    input RXPOLARITY;
    input RXRESET;
    input RXSLIDE;
    input RXUSRCLK2;
    input RXUSRCLK;
    input TSTCLK0;
    input TSTCLK1;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDLYALIGNDISABLE;
    input TXDLYALIGNMONENB;
    input TXDLYALIGNOVERRIDE;
    input TXDLYALIGNRESET;
    input TXDLYALIGNUPDSW;
    input TXELECIDLE;
    input TXENC8B10BUSE;
    input TXENPMAPHASEALIGN;
    input TXINHIBIT;
    input TXPDOWNASYNCH;
    input TXPLLLKDETEN;
    input TXPLLPOWERDOWN;
    input TXPMASETPHASE;
    input TXPOLARITY;
    input TXPRBSFORCEERR;
    input TXRESET;
    input TXSTARTSEQ;
    input TXSWING;
    input TXUSRCLK2;
    input TXUSRCLK;
    input USRCODEERR;
    input [12:0] GTXTEST;
    input [15:0] DI;
    input [19:0] TSTIN;
    input [1:0] MGTREFCLKRX;
    input [1:0] MGTREFCLKTX;
    input [1:0] NORTHREFCLKRX;
    input [1:0] NORTHREFCLKTX;
    input [1:0] RXPOWERDOWN;
    input [1:0] RXRATE;
    input [1:0] SOUTHREFCLKRX;
    input [1:0] SOUTHREFCLKTX;
    input [1:0] TXPOWERDOWN;
    input [1:0] TXRATE;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXENPRBSTST;
    input [2:0] RXPLLREFSELDY;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXENPRBSTST;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXPLLREFSELDY;
    input [31:0] TXDATA;
    input [3:0] DFETAP3;
    input [3:0] DFETAP4;
    input [3:0] RXCHBONDI;
    input [3:0] TXBYPASS8B10B;
    input [3:0] TXCHARDISPMODE;
    input [3:0] TXCHARDISPVAL;
    input [3:0] TXCHARISK;
    input [3:0] TXDIFFCTRL;
    input [3:0] TXPREEMPHASIS;
    input [4:0] DFETAP1;
    input [4:0] DFETAP2;
    input [4:0] TXPOSTEMPHASIS;
    input [5:0] DFECLKDLYADJ;
    input [6:0] TXSEQUENCE;
    input [7:0] DADDR;
    input [9:0] RXEQMIX;
endmodule

module IBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IFD_DELAY_VALUE = "AUTO";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDS_GTHE1 (...);
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFG (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
endmodule

module IBUFGDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter DIFF_TERM = "FALSE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFGDS_DIFF_OUT (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    output OB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

(* keep *)
module IDELAYCTRL (...);
    parameter SIM_DEVICE = "7SERIES";
    output RDY;
    (* clkbuf_sink *)
    input REFCLK;
    input RST;
endmodule

module IOBUF (...);
    parameter integer DRIVE = 12;
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    output O;
    (* iopad_external_pin *)
    inout IO;
    input I;
    input T;
endmodule

module IOBUFDS (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    output O;
    (* iopad_external_pin *)
    inout IO;
    inout IOB;
    input I;
    input T;
endmodule

module IODELAYE1 (...);
    parameter CINVCTRL_SEL = "FALSE";
    parameter DELAY_SRC = "I";
    parameter HIGH_PERFORMANCE_MODE = "FALSE";
    parameter IDELAY_TYPE = "DEFAULT";
    parameter integer IDELAY_VALUE = 0;
    parameter ODELAY_TYPE = "FIXED";
    parameter integer ODELAY_VALUE = 0;
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    output [4:0] CNTVALUEOUT;
    output DATAOUT;
    (* clkbuf_sink *)
    input C;
    input CE;
    input CINVCTRL;
    input CLKIN;
    input [4:0] CNTVALUEIN;
    input DATAIN;
    input IDATAIN;
    input INC;
    input ODATAIN;
    input RST;
    input T;
endmodule

module ISERDESE1 (...);
    parameter DATA_RATE = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter DYN_CLKDIV_INV_EN = "FALSE";
    parameter DYN_CLK_INV_EN = "FALSE";
    parameter [0:0] INIT_Q1 = 1'b0;
    parameter [0:0] INIT_Q2 = 1'b0;
    parameter [0:0] INIT_Q3 = 1'b0;
    parameter [0:0] INIT_Q4 = 1'b0;
    parameter INTERFACE_TYPE = "MEMORY";
    parameter integer NUM_CE = 2;
    parameter IOBDELAY = "NONE";
    parameter OFB_USED = "FALSE";
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_Q1 = 1'b0;
    parameter [0:0] SRVAL_Q2 = 1'b0;
    parameter [0:0] SRVAL_Q3 = 1'b0;
    parameter [0:0] SRVAL_Q4 = 1'b0;
    output O;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output SHIFTOUT1;
    output SHIFTOUT2;
    input BITSLIP;
    input CE1;
    input CE2;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKB;
    (* clkbuf_sink *)
    input CLKDIV;
    input D;
    input DDLY;
    input DYNCLKDIVSEL;
    input DYNCLKSEL;
    (* clkbuf_sink *)
    input OCLK;
    input OFB;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
endmodule

module KEEPER (...);
    inout O;
endmodule

module OBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
endmodule

module OBUFT (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter integer DRIVE = 12;
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    input I;
    input T;
endmodule

module OBUFTDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
    input T;
endmodule

module OSERDESE1 (...);
    parameter DATA_RATE_OQ = "DDR";
    parameter DATA_RATE_TQ = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter integer DDR3_DATA = 1;
    parameter [0:0] INIT_OQ = 1'b0;
    parameter [0:0] INIT_TQ = 1'b0;
    parameter INTERFACE_TYPE = "DEFAULT";
    parameter integer ODELAY_USED = 0;
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_OQ = 1'b0;
    parameter [0:0] SRVAL_TQ = 1'b0;
    parameter integer TRISTATE_WIDTH = 4;
    output OCBEXTEND;
    output OFB;
    output OQ;
    output SHIFTOUT1;
    output SHIFTOUT2;
    output TFB;
    output TQ;
    (* clkbuf_sink *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    input CLKPERF;
    input CLKPERFDELAY;
    input D1;
    input D2;
    input D3;
    input D4;
    input D5;
    input D6;
    input OCE;
    input ODV;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
    input T1;
    input T2;
    input T3;
    input T4;
    input TCE;
    input WC;
endmodule

module PULLDOWN (...);
    output O;
endmodule

module PULLUP (...);
    output O;
endmodule

module TEMAC_SINGLE (...);
    parameter EMAC_1000BASEX_ENABLE = "FALSE";
    parameter EMAC_ADDRFILTER_ENABLE = "FALSE";
    parameter EMAC_BYTEPHY = "FALSE";
    parameter EMAC_CTRLLENCHECK_DISABLE = "FALSE";
    parameter [0:7] EMAC_DCRBASEADDR = 8'h00;
    parameter EMAC_GTLOOPBACK = "FALSE";
    parameter EMAC_HOST_ENABLE = "FALSE";
    parameter [8:0] EMAC_LINKTIMERVAL = 9'h000;
    parameter EMAC_LTCHECK_DISABLE = "FALSE";
    parameter EMAC_MDIO_ENABLE = "FALSE";
    parameter EMAC_MDIO_IGNORE_PHYADZERO = "FALSE";
    parameter [47:0] EMAC_PAUSEADDR = 48'h000000000000;
    parameter EMAC_PHYINITAUTONEG_ENABLE = "FALSE";
    parameter EMAC_PHYISOLATE = "FALSE";
    parameter EMAC_PHYLOOPBACKMSB = "FALSE";
    parameter EMAC_PHYPOWERDOWN = "FALSE";
    parameter EMAC_PHYRESET = "FALSE";
    parameter EMAC_RGMII_ENABLE = "FALSE";
    parameter EMAC_RX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC_RXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC_RXHALFDUPLEX = "FALSE";
    parameter EMAC_RXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC_RXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC_RXRESET = "FALSE";
    parameter EMAC_RXVLAN_ENABLE = "FALSE";
    parameter EMAC_RX_ENABLE = "TRUE";
    parameter EMAC_SGMII_ENABLE = "FALSE";
    parameter EMAC_SPEED_LSB = "FALSE";
    parameter EMAC_SPEED_MSB = "FALSE";
    parameter EMAC_TX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC_TXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC_TXHALFDUPLEX = "FALSE";
    parameter EMAC_TXIFGADJUST_ENABLE = "FALSE";
    parameter EMAC_TXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC_TXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC_TXRESET = "FALSE";
    parameter EMAC_TXVLAN_ENABLE = "FALSE";
    parameter EMAC_TX_ENABLE = "TRUE";
    parameter [47:0] EMAC_UNICASTADDR = 48'h000000000000;
    parameter EMAC_UNIDIRECTION_ENABLE = "FALSE";
    parameter EMAC_USECLKEN = "FALSE";
    parameter SIM_VERSION = "1.0";
    output DCRHOSTDONEIR;
    output EMACCLIENTANINTERRUPT;
    output EMACCLIENTRXBADFRAME;
    output EMACCLIENTRXCLIENTCLKOUT;
    output EMACCLIENTRXDVLD;
    output EMACCLIENTRXDVLDMSW;
    output EMACCLIENTRXFRAMEDROP;
    output EMACCLIENTRXGOODFRAME;
    output EMACCLIENTRXSTATSBYTEVLD;
    output EMACCLIENTRXSTATSVLD;
    output EMACCLIENTTXACK;
    output EMACCLIENTTXCLIENTCLKOUT;
    output EMACCLIENTTXCOLLISION;
    output EMACCLIENTTXRETRANSMIT;
    output EMACCLIENTTXSTATS;
    output EMACCLIENTTXSTATSBYTEVLD;
    output EMACCLIENTTXSTATSVLD;
    output EMACDCRACK;
    output EMACPHYENCOMMAALIGN;
    output EMACPHYLOOPBACKMSB;
    output EMACPHYMCLKOUT;
    output EMACPHYMDOUT;
    output EMACPHYMDTRI;
    output EMACPHYMGTRXRESET;
    output EMACPHYMGTTXRESET;
    output EMACPHYPOWERDOWN;
    output EMACPHYSYNCACQSTATUS;
    output EMACPHYTXCHARDISPMODE;
    output EMACPHYTXCHARDISPVAL;
    output EMACPHYTXCHARISK;
    output EMACPHYTXCLK;
    output EMACPHYTXEN;
    output EMACPHYTXER;
    output EMACPHYTXGMIIMIICLKOUT;
    output EMACSPEEDIS10100;
    output HOSTMIIMRDY;
    output [0:31] EMACDCRDBUS;
    output [15:0] EMACCLIENTRXD;
    output [31:0] HOSTRDDATA;
    output [6:0] EMACCLIENTRXSTATS;
    output [7:0] EMACPHYTXD;
    input CLIENTEMACDCMLOCKED;
    input CLIENTEMACPAUSEREQ;
    input CLIENTEMACRXCLIENTCLKIN;
    input CLIENTEMACTXCLIENTCLKIN;
    input CLIENTEMACTXDVLD;
    input CLIENTEMACTXDVLDMSW;
    input CLIENTEMACTXFIRSTBYTE;
    input CLIENTEMACTXUNDERRUN;
    input DCREMACCLK;
    input DCREMACENABLE;
    input DCREMACREAD;
    input DCREMACWRITE;
    input HOSTCLK;
    input HOSTMIIMSEL;
    input HOSTREQ;
    input PHYEMACCOL;
    input PHYEMACCRS;
    input PHYEMACGTXCLK;
    input PHYEMACMCLKIN;
    input PHYEMACMDIN;
    input PHYEMACMIITXCLK;
    input PHYEMACRXCHARISCOMMA;
    input PHYEMACRXCHARISK;
    input PHYEMACRXCLK;
    input PHYEMACRXDISPERR;
    input PHYEMACRXDV;
    input PHYEMACRXER;
    input PHYEMACRXNOTINTABLE;
    input PHYEMACRXRUNDISP;
    input PHYEMACSIGNALDET;
    input PHYEMACTXBUFERR;
    input PHYEMACTXGMIIMIICLKIN;
    input RESET;
    input [0:31] DCREMACDBUS;
    input [0:9] DCREMACABUS;
    input [15:0] CLIENTEMACPAUSEVAL;
    input [15:0] CLIENTEMACTXD;
    input [1:0] HOSTOPCODE;
    input [1:0] PHYEMACRXBUFSTATUS;
    input [2:0] PHYEMACRXCLKCORCNT;
    input [31:0] HOSTWRDATA;
    input [4:0] PHYEMACPHYAD;
    input [7:0] CLIENTEMACTXIFGDELAY;
    input [7:0] PHYEMACRXD;
    input [9:0] HOSTADDR;
endmodule

module FIFO18E1 (...);
    parameter ALMOST_EMPTY_OFFSET = 13'h0080;
    parameter ALMOST_FULL_OFFSET = 13'h0080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_SYN = "FALSE";
    parameter FIFO_MODE = "FIFO18";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter INIT = 36'h0;
    parameter SIM_DEVICE = "VIRTEX6";
    parameter SRVAL = 36'h0;
    parameter IS_RDCLK_INVERTED = 1'b0;
    parameter IS_RDEN_INVERTED = 1'b0;
    parameter IS_RSTREG_INVERTED = 1'b0;
    parameter IS_RST_INVERTED = 1'b0;
    parameter IS_WRCLK_INVERTED = 1'b0;
    parameter IS_WREN_INVERTED = 1'b0;
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [31:0] DO;
    output [3:0] DOP;
    output EMPTY;
    output FULL;
    output [11:0] RDCOUNT;
    output RDERR;
    output [11:0] WRCOUNT;
    output WRERR;
    input [31:0] DI;
    input [3:0] DIP;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input REGCE;
    input RST;
    input RSTREG;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module FIFO36E1 (...);
    parameter ALMOST_EMPTY_OFFSET = 13'h0080;
    parameter ALMOST_FULL_OFFSET = 13'h0080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter EN_SYN = "FALSE";
    parameter FIFO_MODE = "FIFO36";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter INIT = 72'h0;
    parameter SIM_DEVICE = "VIRTEX6";
    parameter SRVAL = 72'h0;
    parameter IS_RDCLK_INVERTED = 1'b0;
    parameter IS_RDEN_INVERTED = 1'b0;
    parameter IS_RSTREG_INVERTED = 1'b0;
    parameter IS_RST_INVERTED = 1'b0;
    parameter IS_WRCLK_INVERTED = 1'b0;
    parameter IS_WREN_INVERTED = 1'b0;
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output DBITERR;
    output [63:0] DO;
    output [7:0] DOP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output SBITERR;
    output [12:0] WRCOUNT;
    output WRERR;
    input [63:0] DI;
    input [7:0] DIP;
    input INJECTDBITERR;
    input INJECTSBITERR;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input REGCE;
    input RST;
    input RSTREG;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
endmodule

module RAM128X1S (...);
    parameter [127:0] INIT = 128'h00000000000000000000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input A6;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM256X1S (...);
    parameter [255:0] INIT = 256'h0;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input [7:0] A;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32M (...);
    parameter [63:0] INIT_A = 64'h0000000000000000;
    parameter [63:0] INIT_B = 64'h0000000000000000;
    parameter [63:0] INIT_C = 64'h0000000000000000;
    parameter [63:0] INIT_D = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output [1:0] DOA;
    output [1:0] DOB;
    output [1:0] DOC;
    output [1:0] DOD;
    input [4:0] ADDRA;
    input [4:0] ADDRB;
    input [4:0] ADDRC;
    input [4:0] ADDRD;
    input [1:0] DIA;
    input [1:0] DIB;
    input [1:0] DIC;
    input [1:0] DID;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32X1S (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32X1S_1 (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM32X2S (...);
    parameter [31:0] INIT_00 = 32'h00000000;
    parameter [31:0] INIT_01 = 32'h00000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O0;
    output O1;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input D0;
    input D1;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64M (...);
    parameter [63:0] INIT_A = 64'h0000000000000000;
    parameter [63:0] INIT_B = 64'h0000000000000000;
    parameter [63:0] INIT_C = 64'h0000000000000000;
    parameter [63:0] INIT_D = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output DOA;
    output DOB;
    output DOC;
    output DOD;
    input [5:0] ADDRA;
    input [5:0] ADDRB;
    input [5:0] ADDRC;
    input [5:0] ADDRD;
    input DIA;
    input DIB;
    input DIC;
    input DID;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64X1S (...);
    parameter [63:0] INIT = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64X1S_1 (...);
    parameter [63:0] INIT = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input D;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module RAM64X2S (...);
    parameter [63:0] INIT_00 = 64'h0000000000000000;
    parameter [63:0] INIT_01 = 64'h0000000000000000;
    parameter [0:0] IS_WCLK_INVERTED = 1'b0;
    output O0;
    output O1;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input D0;
    input D1;
    (* clkbuf_sink *)
    input WCLK;
    input WE;
endmodule

module ROM128X1 (...);
    parameter [127:0] INIT = 128'h00000000000000000000000000000000;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input A6;
endmodule

module ROM256X1 (...);
    parameter [255:0] INIT = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
    input A6;
    input A7;
endmodule

module ROM32X1 (...);
    parameter [31:0] INIT = 32'h00000000;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
endmodule

module ROM64X1 (...);
    parameter [63:0] INIT = 64'h0000000000000000;
    output O;
    input A0;
    input A1;
    input A2;
    input A3;
    input A4;
    input A5;
endmodule

module IDDR (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter INIT_Q1 = 1'b0;
    parameter INIT_Q2 = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter SRTYPE = "SYNC";
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    input C;
    input CE;
    input D;
    input R;
    input S;
endmodule

module IDDR_2CLK (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter INIT_Q1 = 1'b0;
    parameter INIT_Q2 = 1'b0;
    parameter [0:0] IS_CB_INVERTED = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter SRTYPE = "SYNC";
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    input C;
    (* clkbuf_sink *)
    input CB;
    input CE;
    input D;
    input R;
    input S;
endmodule

module LDCE (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_G_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    input CLR;
    input D;
    input G;
    input GE;
endmodule

module LDPE (...);
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_G_INVERTED = 1'b0;
    parameter [0:0] IS_PRE_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    input D;
    input G;
    input GE;
    input PRE;
endmodule

module ODDR (...);
    output Q;
    (* clkbuf_sink *)
    input C;
    input CE;
    input D1;
    input D2;
    input R;
    input S;
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter INIT = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter SRTYPE = "SYNC";
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
endmodule

module CFGLUT5 (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    output CDO;
    output O5;
    output O6;
    input I4;
    input I3;
    input I2;
    input I1;
    input I0;
    input CDI;
    input CE;
    (* clkbuf_sink *)
    input CLK;
endmodule

