// Flip-flop D
module  \$_DFF_P_ (input D, input C, output Q);
   parameter WYSIWYG="TRUE";
   dffeas #(.is_wysiwyg(WYSIWYG)) _TECHMAP_REPLACE_ (.d(D), .q(Q), .clk(C), .clrn(1'b1), .prn(1'b1), .ena(1'b1), .asdata(1'b0), .aload(1'b0), .sclr(1'b0), .sload(1'b0));
endmodule //

// Input buffer map
module \$__inpad (input I, output O);
    cycloneiv_io_ibuf _TECHMAP_REPLACE_ (.o(O), .i(I), .ibar(1'b0));
endmodule 

// Output buffer map   
module \$__outpad (input I, output O);
    cycloneiv_io_obuf _TECHMAP_REPLACE_ (.o(O), .i(I), .oe(1'b1));
endmodule 

// LUT Map
/* 0 -> datac
   1 -> cin */
module \$lut (A, Y);
   parameter WIDTH  = 0;
   parameter LUT    = 0;
   parameter SPLIT4 = {LUT[15:12], LUT[7:4], LUT[11:8], LUT[3:0]}; // used for 4-in luts, KISS;
   input [WIDTH-1:0] A;
   output 	     Y;
   generate 
      if (WIDTH == 1) begin
	   assign Y = ~A[0]; // Not need to spend 1 logic cell for such an easy function
      end else
      if (WIDTH == 2) begin
           cycloneiv_lcell_comb #(.lut_mask({4{LUT}}), .sum_lutc_input("datac")) _TECHMAP_REPLACE_ (.combout(Y), .dataa(A[0]), .datab(A[1]), .datac(1'b1),.datad(1'b1));
      end else
      if(WIDTH == 3) begin 
	   cycloneiv_lcell_comb #(.lut_mask({2{LUT}}), .sum_lutc_input("datac")) _TECHMAP_REPLACE_ (.combout(Y), .dataa(A[0]), .datab(A[1]), .datac(A[2]),.datad(1'b1));
      end else
      if(WIDTH == 4) begin
	   cycloneiv_lcell_comb #(.lut_mask(LUT), .sum_lutc_input("datac")) _TECHMAP_REPLACE_ (.combout(Y), .dataa(A[0]), .datab(A[1]), .datac(A[2]),.datad(A[3]));
      end else
	   wire _TECHMAP_FAIL_ = 1;
   endgenerate
endmodule //

	    
