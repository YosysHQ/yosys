`define parvez ahmad
`define  WIRE wire
`define TEN 10

module `parvez();
parameter param = `TEN;
`WIRE w;
assign w = `TEN;
endmodule
