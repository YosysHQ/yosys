module adder(sum , co, a, b, ci);
output	reg		[31:0]	sum;
output	reg				co;
input	wire	[31:0]	a, b;
input wire				ci;
endmodule
