module test(input in, output out);
assign out = 1'b1;
endmodule
