module a;
wire [5:0]x;
wire [3:0]y;
assign y = x 55;
endmodule

