module test(A, B, Y);
    input  [1:0] A, B;
    output [1:0] Y = A * B;
endmodule
