`default_nettype none
module latch_1990_gate
  (output wire [1:0] x);
   assign x = 2'b10;
endmodule // latch_1990_gate

