module my_module(
    input a,
    input b,
    output y
);
   // Perform operation
   assign y = a | b;

endmodule
